/*  
Copyright 2019 XCrypt Studio                
																	 
Licensed under the Apache License, Version 2.0 (the "License");         
you may not use this file except in compliance with the License.        
You may obtain a copy of the License at                                 
																	 
 http://www.apache.org/licenses/LICENSE-2.0                          
																	 
Unless required by applicable law or agreed to in writing, software    
distributed under the License is distributed on an "AS IS" BASIS,       
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and     
limitations under the License.                                          
*/  

// ------------------------------------------------------------------------------
// File name        :   cast5_sbox3.v
// Function         :   CAST5 Cryptographic Algorithm Core SBox-3 & SBox-7
// ------------------------------------------------------------------------------
// Author           :   Xie
// Version          ：  v-1.0
// Date				:   2019-2-2
// Email            :   xcrypt@126.com
// ------------------------------------------------------------------------------

`timescale 1ns / 1ps

module cast5_sbox37(
	input 			i_clk,
	input			i_sel, //1:s-box3 0:s-box7
    input   [7:0]   i_addr,
    output  [31:0]  o_data
    );
	
	localparam DLY = 1;
	
    reg [31:0] r_dout;
    assign o_data = r_dout;
	//
    always@(posedge i_clk) begin
		if(i_sel) begin		//sbox-3
			case(i_addr)
				8'h00 : r_dout <= #DLY 32'h8defc240;
				8'h01 : r_dout <= #DLY 32'h25fa5d9f;
				8'h02 : r_dout <= #DLY 32'heb903dbf;
				8'h03 : r_dout <= #DLY 32'he810c907;
				8'h04 : r_dout <= #DLY 32'h47607fff;
				8'h05 : r_dout <= #DLY 32'h369fe44b;
				8'h06 : r_dout <= #DLY 32'h8c1fc644;
				8'h07 : r_dout <= #DLY 32'haececa90;
				8'h08 : r_dout <= #DLY 32'hbeb1f9bf;
				8'h09 : r_dout <= #DLY 32'heefbcaea;
				8'h0a : r_dout <= #DLY 32'he8cf1950;
				8'h0b : r_dout <= #DLY 32'h51df07ae;
				8'h0c : r_dout <= #DLY 32'h920e8806;
				8'h0d : r_dout <= #DLY 32'hf0ad0548;
				8'h0e : r_dout <= #DLY 32'he13c8d83;
				8'h0f : r_dout <= #DLY 32'h927010d5;
				8'h10 : r_dout <= #DLY 32'h11107d9f;
				8'h11 : r_dout <= #DLY 32'h07647db9;
				8'h12 : r_dout <= #DLY 32'hb2e3e4d4;
				8'h13 : r_dout <= #DLY 32'h3d4f285e;
				8'h14 : r_dout <= #DLY 32'hb9afa820;
				8'h15 : r_dout <= #DLY 32'hfade82e0;
				8'h16 : r_dout <= #DLY 32'ha067268b;
				8'h17 : r_dout <= #DLY 32'h8272792e;
				8'h18 : r_dout <= #DLY 32'h553fb2c0;
				8'h19 : r_dout <= #DLY 32'h489ae22b;
				8'h1a : r_dout <= #DLY 32'hd4ef9794;
				8'h1b : r_dout <= #DLY 32'h125e3fbc;
				8'h1c : r_dout <= #DLY 32'h21fffcee;
				8'h1d : r_dout <= #DLY 32'h825b1bfd;
				8'h1e : r_dout <= #DLY 32'h9255c5ed;
				8'h1f : r_dout <= #DLY 32'h1257a240;
				8'h20 : r_dout <= #DLY 32'h4e1a8302;
				8'h21 : r_dout <= #DLY 32'hbae07fff;
				8'h22 : r_dout <= #DLY 32'h528246e7;
				8'h23 : r_dout <= #DLY 32'h8e57140e;
				8'h24 : r_dout <= #DLY 32'h3373f7bf;
				8'h25 : r_dout <= #DLY 32'h8c9f8188;
				8'h26 : r_dout <= #DLY 32'ha6fc4ee8;
				8'h27 : r_dout <= #DLY 32'hc982b5a5;
				8'h28 : r_dout <= #DLY 32'ha8c01db7;
				8'h29 : r_dout <= #DLY 32'h579fc264;
				8'h2a : r_dout <= #DLY 32'h67094f31;
				8'h2b : r_dout <= #DLY 32'hf2bd3f5f;
				8'h2c : r_dout <= #DLY 32'h40fff7c1;
				8'h2d : r_dout <= #DLY 32'h1fb78dfc;
				8'h2e : r_dout <= #DLY 32'h8e6bd2c1;
				8'h2f : r_dout <= #DLY 32'h437be59b;
				8'h30 : r_dout <= #DLY 32'h99b03dbf;
				8'h31 : r_dout <= #DLY 32'hb5dbc64b;
				8'h32 : r_dout <= #DLY 32'h638dc0e6;
				8'h33 : r_dout <= #DLY 32'h55819d99;
				8'h34 : r_dout <= #DLY 32'ha197c81c;
				8'h35 : r_dout <= #DLY 32'h4a012d6e;
				8'h36 : r_dout <= #DLY 32'hc5884a28;
				8'h37 : r_dout <= #DLY 32'hccc36f71;
				8'h38 : r_dout <= #DLY 32'hb843c213;
				8'h39 : r_dout <= #DLY 32'h6c0743f1;
				8'h3a : r_dout <= #DLY 32'h8309893c;
				8'h3b : r_dout <= #DLY 32'h0feddd5f;
				8'h3c : r_dout <= #DLY 32'h2f7fe850;
				8'h3d : r_dout <= #DLY 32'hd7c07f7e;
				8'h3e : r_dout <= #DLY 32'h02507fbf;
				8'h3f : r_dout <= #DLY 32'h5afb9a04;
				8'h40 : r_dout <= #DLY 32'ha747d2d0;
				8'h41 : r_dout <= #DLY 32'h1651192e;
				8'h42 : r_dout <= #DLY 32'haf70bf3e;
				8'h43 : r_dout <= #DLY 32'h58c31380;
				8'h44 : r_dout <= #DLY 32'h5f98302e;
				8'h45 : r_dout <= #DLY 32'h727cc3c4;
				8'h46 : r_dout <= #DLY 32'h0a0fb402;
				8'h47 : r_dout <= #DLY 32'h0f7fef82;
				8'h48 : r_dout <= #DLY 32'h8c96fdad;
				8'h49 : r_dout <= #DLY 32'h5d2c2aae;
				8'h4a : r_dout <= #DLY 32'h8ee99a49;
				8'h4b : r_dout <= #DLY 32'h50da88b8;
				8'h4c : r_dout <= #DLY 32'h8427f4a0;
				8'h4d : r_dout <= #DLY 32'h1eac5790;
				8'h4e : r_dout <= #DLY 32'h796fb449;
				8'h4f : r_dout <= #DLY 32'h8252dc15;
				8'h50 : r_dout <= #DLY 32'hefbd7d9b;
				8'h51 : r_dout <= #DLY 32'ha672597d;
				8'h52 : r_dout <= #DLY 32'hada840d8;
				8'h53 : r_dout <= #DLY 32'h45f54504;
				8'h54 : r_dout <= #DLY 32'hfa5d7403;
				8'h55 : r_dout <= #DLY 32'he83ec305;
				8'h56 : r_dout <= #DLY 32'h4f91751a;
				8'h57 : r_dout <= #DLY 32'h925669c2;
				8'h58 : r_dout <= #DLY 32'h23efe941;
				8'h59 : r_dout <= #DLY 32'ha903f12e;
				8'h5a : r_dout <= #DLY 32'h60270df2;
				8'h5b : r_dout <= #DLY 32'h0276e4b6;
				8'h5c : r_dout <= #DLY 32'h94fd6574;
				8'h5d : r_dout <= #DLY 32'h927985b2;
				8'h5e : r_dout <= #DLY 32'h8276dbcb;
				8'h5f : r_dout <= #DLY 32'h02778176;
				8'h60 : r_dout <= #DLY 32'hf8af918d;
				8'h61 : r_dout <= #DLY 32'h4e48f79e;
				8'h62 : r_dout <= #DLY 32'h8f616ddf;
				8'h63 : r_dout <= #DLY 32'he29d840e;
				8'h64 : r_dout <= #DLY 32'h842f7d83;
				8'h65 : r_dout <= #DLY 32'h340ce5c8;
				8'h66 : r_dout <= #DLY 32'h96bbb682;
				8'h67 : r_dout <= #DLY 32'h93b4b148;
				8'h68 : r_dout <= #DLY 32'hef303cab;
				8'h69 : r_dout <= #DLY 32'h984faf28;
				8'h6a : r_dout <= #DLY 32'h779faf9b;
				8'h6b : r_dout <= #DLY 32'h92dc560d;
				8'h6c : r_dout <= #DLY 32'h224d1e20;
				8'h6d : r_dout <= #DLY 32'h8437aa88;
				8'h6e : r_dout <= #DLY 32'h7d29dc96;
				8'h6f : r_dout <= #DLY 32'h2756d3dc;
				8'h70 : r_dout <= #DLY 32'h8b907cee;
				8'h71 : r_dout <= #DLY 32'hb51fd240;
				8'h72 : r_dout <= #DLY 32'he7c07ce3;
				8'h73 : r_dout <= #DLY 32'he566b4a1;
				8'h74 : r_dout <= #DLY 32'hc3e9615e;
				8'h75 : r_dout <= #DLY 32'h3cf8209d;
				8'h76 : r_dout <= #DLY 32'h6094d1e3;
				8'h77 : r_dout <= #DLY 32'hcd9ca341;
				8'h78 : r_dout <= #DLY 32'h5c76460e;
				8'h79 : r_dout <= #DLY 32'h00ea983b;
				8'h7a : r_dout <= #DLY 32'hd4d67881;
				8'h7b : r_dout <= #DLY 32'hfd47572c;
				8'h7c : r_dout <= #DLY 32'hf76cedd9;
				8'h7d : r_dout <= #DLY 32'hbda8229c;
				8'h7e : r_dout <= #DLY 32'h127dadaa;
				8'h7f : r_dout <= #DLY 32'h438a074e;
				8'h80 : r_dout <= #DLY 32'h1f97c090;
				8'h81 : r_dout <= #DLY 32'h081bdb8a;
				8'h82 : r_dout <= #DLY 32'h93a07ebe;
				8'h83 : r_dout <= #DLY 32'hb938ca15;
				8'h84 : r_dout <= #DLY 32'h97b03cff;
				8'h85 : r_dout <= #DLY 32'h3dc2c0f8;
				8'h86 : r_dout <= #DLY 32'h8d1ab2ec;
				8'h87 : r_dout <= #DLY 32'h64380e51;
				8'h88 : r_dout <= #DLY 32'h68cc7bfb;
				8'h89 : r_dout <= #DLY 32'hd90f2788;
				8'h8a : r_dout <= #DLY 32'h12490181;
				8'h8b : r_dout <= #DLY 32'h5de5ffd4;
				8'h8c : r_dout <= #DLY 32'hdd7ef86a;
				8'h8d : r_dout <= #DLY 32'h76a2e214;
				8'h8e : r_dout <= #DLY 32'hb9a40368;
				8'h8f : r_dout <= #DLY 32'h925d958f;
				8'h90 : r_dout <= #DLY 32'h4b39fffa;
				8'h91 : r_dout <= #DLY 32'hba39aee9;
				8'h92 : r_dout <= #DLY 32'ha4ffd30b;
				8'h93 : r_dout <= #DLY 32'hfaf7933b;
				8'h94 : r_dout <= #DLY 32'h6d498623;
				8'h95 : r_dout <= #DLY 32'h193cbcfa;
				8'h96 : r_dout <= #DLY 32'h27627545;
				8'h97 : r_dout <= #DLY 32'h825cf47a;
				8'h98 : r_dout <= #DLY 32'h61bd8ba0;
				8'h99 : r_dout <= #DLY 32'hd11e42d1;
				8'h9a : r_dout <= #DLY 32'hcead04f4;
				8'h9b : r_dout <= #DLY 32'h127ea392;
				8'h9c : r_dout <= #DLY 32'h10428db7;
				8'h9d : r_dout <= #DLY 32'h8272a972;
				8'h9e : r_dout <= #DLY 32'h9270c4a8;
				8'h9f : r_dout <= #DLY 32'h127de50b;
				8'ha0 : r_dout <= #DLY 32'h285ba1c8;
				8'ha1 : r_dout <= #DLY 32'h3c62f44f;
				8'ha2 : r_dout <= #DLY 32'h35c0eaa5;
				8'ha3 : r_dout <= #DLY 32'he805d231;
				8'ha4 : r_dout <= #DLY 32'h428929fb;
				8'ha5 : r_dout <= #DLY 32'hb4fcdf82;
				8'ha6 : r_dout <= #DLY 32'h4fb66a53;
				8'ha7 : r_dout <= #DLY 32'h0e7dc15b;
				8'ha8 : r_dout <= #DLY 32'h1f081fab;
				8'ha9 : r_dout <= #DLY 32'h108618ae;
				8'haa : r_dout <= #DLY 32'hfcfd086d;
				8'hab : r_dout <= #DLY 32'hf9ff2889;
				8'hac : r_dout <= #DLY 32'h694bcc11;
				8'had : r_dout <= #DLY 32'h236a5cae;
				8'hae : r_dout <= #DLY 32'h12deca4d;
				8'haf : r_dout <= #DLY 32'h2c3f8cc5;
				8'hb0 : r_dout <= #DLY 32'hd2d02dfe;
				8'hb1 : r_dout <= #DLY 32'hf8ef5896;
				8'hb2 : r_dout <= #DLY 32'he4cf52da;
				8'hb3 : r_dout <= #DLY 32'h95155b67;
				8'hb4 : r_dout <= #DLY 32'h494a488c;
				8'hb5 : r_dout <= #DLY 32'hb9b6a80c;
				8'hb6 : r_dout <= #DLY 32'h5c8f82bc;
				8'hb7 : r_dout <= #DLY 32'h89d36b45;
				8'hb8 : r_dout <= #DLY 32'h3a609437;
				8'hb9 : r_dout <= #DLY 32'hec00c9a9;
				8'hba : r_dout <= #DLY 32'h44715253;
				8'hbb : r_dout <= #DLY 32'h0a874b49;
				8'hbc : r_dout <= #DLY 32'hd773bc40;
				8'hbd : r_dout <= #DLY 32'h7c34671c;
				8'hbe : r_dout <= #DLY 32'h02717ef6;
				8'hbf : r_dout <= #DLY 32'h4feb5536;
				8'hc0 : r_dout <= #DLY 32'ha2d02fff;
				8'hc1 : r_dout <= #DLY 32'hd2bf60c4;
				8'hc2 : r_dout <= #DLY 32'hd43f03c0;
				8'hc3 : r_dout <= #DLY 32'h50b4ef6d;
				8'hc4 : r_dout <= #DLY 32'h07478cd1;
				8'hc5 : r_dout <= #DLY 32'h006e1888;
				8'hc6 : r_dout <= #DLY 32'ha2e53f55;
				8'hc7 : r_dout <= #DLY 32'hb9e6d4bc;
				8'hc8 : r_dout <= #DLY 32'ha2048016;
				8'hc9 : r_dout <= #DLY 32'h97573833;
				8'hca : r_dout <= #DLY 32'hd7207d67;
				8'hcb : r_dout <= #DLY 32'hde0f8f3d;
				8'hcc : r_dout <= #DLY 32'h72f87b33;
				8'hcd : r_dout <= #DLY 32'habcc4f33;
				8'hce : r_dout <= #DLY 32'h7688c55d;
				8'hcf : r_dout <= #DLY 32'h7b00a6b0;
				8'hd0 : r_dout <= #DLY 32'h947b0001;
				8'hd1 : r_dout <= #DLY 32'h570075d2;
				8'hd2 : r_dout <= #DLY 32'hf9bb88f8;
				8'hd3 : r_dout <= #DLY 32'h8942019e;
				8'hd4 : r_dout <= #DLY 32'h4264a5ff;
				8'hd5 : r_dout <= #DLY 32'h856302e0;
				8'hd6 : r_dout <= #DLY 32'h72dbd92b;
				8'hd7 : r_dout <= #DLY 32'hee971b69;
				8'hd8 : r_dout <= #DLY 32'h6ea22fde;
				8'hd9 : r_dout <= #DLY 32'h5f08ae2b;
				8'hda : r_dout <= #DLY 32'haf7a616d;
				8'hdb : r_dout <= #DLY 32'he5c98767;
				8'hdc : r_dout <= #DLY 32'hcf1febd2;
				8'hdd : r_dout <= #DLY 32'h61efc8c2;
				8'hde : r_dout <= #DLY 32'hf1ac2571;
				8'hdf : r_dout <= #DLY 32'hcc8239c2;
				8'he0 : r_dout <= #DLY 32'h67214cb8;
				8'he1 : r_dout <= #DLY 32'hb1e583d1;
				8'he2 : r_dout <= #DLY 32'hb7dc3e62;
				8'he3 : r_dout <= #DLY 32'h7f10bdce;
				8'he4 : r_dout <= #DLY 32'hf90a5c38;
				8'he5 : r_dout <= #DLY 32'h0ff0443d;
				8'he6 : r_dout <= #DLY 32'h606e6dc6;
				8'he7 : r_dout <= #DLY 32'h60543a49;
				8'he8 : r_dout <= #DLY 32'h5727c148;
				8'he9 : r_dout <= #DLY 32'h2be98a1d;
				8'hea : r_dout <= #DLY 32'h8ab41738;
				8'heb : r_dout <= #DLY 32'h20e1be24;
				8'hec : r_dout <= #DLY 32'haf96da0f;
				8'hed : r_dout <= #DLY 32'h68458425;
				8'hee : r_dout <= #DLY 32'h99833be5;
				8'hef : r_dout <= #DLY 32'h600d457d;
				8'hf0 : r_dout <= #DLY 32'h282f9350;
				8'hf1 : r_dout <= #DLY 32'h8334b362;
				8'hf2 : r_dout <= #DLY 32'hd91d1120;
				8'hf3 : r_dout <= #DLY 32'h2b6d8da0;
				8'hf4 : r_dout <= #DLY 32'h642b1e31;
				8'hf5 : r_dout <= #DLY 32'h9c305a00;
				8'hf6 : r_dout <= #DLY 32'h52bce688;
				8'hf7 : r_dout <= #DLY 32'h1b03588a;
				8'hf8 : r_dout <= #DLY 32'hf7baefd5;
				8'hf9 : r_dout <= #DLY 32'h4142ed9c;
				8'hfa : r_dout <= #DLY 32'ha4315c11;
				8'hfb : r_dout <= #DLY 32'h83323ec5;
				8'hfc : r_dout <= #DLY 32'hdfef4636;
				8'hfd : r_dout <= #DLY 32'ha133c501;
				8'hfe : r_dout <= #DLY 32'he9d3531c;
				8'hff : r_dout <= #DLY 32'hee353783;
			endcase
		end else begin
			case(i_addr)	//s-box7
				8'h00 : r_dout <= #DLY 32'h85e04019;
				8'h01 : r_dout <= #DLY 32'h332bf567;
				8'h02 : r_dout <= #DLY 32'h662dbfff;
				8'h03 : r_dout <= #DLY 32'hcfc65693;
				8'h04 : r_dout <= #DLY 32'h2a8d7f6f;
				8'h05 : r_dout <= #DLY 32'hab9bc912;
				8'h06 : r_dout <= #DLY 32'hde6008a1;
				8'h07 : r_dout <= #DLY 32'h2028da1f;
				8'h08 : r_dout <= #DLY 32'h0227bce7;
				8'h09 : r_dout <= #DLY 32'h4d642916;
				8'h0a : r_dout <= #DLY 32'h18fac300;
				8'h0b : r_dout <= #DLY 32'h50f18b82;
				8'h0c : r_dout <= #DLY 32'h2cb2cb11;
				8'h0d : r_dout <= #DLY 32'hb232e75c;
				8'h0e : r_dout <= #DLY 32'h4b3695f2;
				8'h0f : r_dout <= #DLY 32'hb28707de;
				8'h10 : r_dout <= #DLY 32'ha05fbcf6;
				8'h11 : r_dout <= #DLY 32'hcd4181e9;
				8'h12 : r_dout <= #DLY 32'he150210c;
				8'h13 : r_dout <= #DLY 32'he24ef1bd;
				8'h14 : r_dout <= #DLY 32'hb168c381;
				8'h15 : r_dout <= #DLY 32'hfde4e789;
				8'h16 : r_dout <= #DLY 32'h5c79b0d8;
				8'h17 : r_dout <= #DLY 32'h1e8bfd43;
				8'h18 : r_dout <= #DLY 32'h4d495001;
				8'h19 : r_dout <= #DLY 32'h38be4341;
				8'h1a : r_dout <= #DLY 32'h913cee1d;
				8'h1b : r_dout <= #DLY 32'h92a79c3f;
				8'h1c : r_dout <= #DLY 32'h089766be;
				8'h1d : r_dout <= #DLY 32'hbaeeadf4;
				8'h1e : r_dout <= #DLY 32'h1286becf;
				8'h1f : r_dout <= #DLY 32'hb6eacb19;
				8'h20 : r_dout <= #DLY 32'h2660c200;
				8'h21 : r_dout <= #DLY 32'h7565bde4;
				8'h22 : r_dout <= #DLY 32'h64241f7a;
				8'h23 : r_dout <= #DLY 32'h8248dca9;
				8'h24 : r_dout <= #DLY 32'hc3b3ad66;
				8'h25 : r_dout <= #DLY 32'h28136086;
				8'h26 : r_dout <= #DLY 32'h0bd8dfa8;
				8'h27 : r_dout <= #DLY 32'h356d1cf2;
				8'h28 : r_dout <= #DLY 32'h107789be;
				8'h29 : r_dout <= #DLY 32'hb3b2e9ce;
				8'h2a : r_dout <= #DLY 32'h0502aa8f;
				8'h2b : r_dout <= #DLY 32'h0bc0351e;
				8'h2c : r_dout <= #DLY 32'h166bf52a;
				8'h2d : r_dout <= #DLY 32'heb12ff82;
				8'h2e : r_dout <= #DLY 32'he3486911;
				8'h2f : r_dout <= #DLY 32'hd34d7516;
				8'h30 : r_dout <= #DLY 32'h4e7b3aff;
				8'h31 : r_dout <= #DLY 32'h5f43671b;
				8'h32 : r_dout <= #DLY 32'h9cf6e037;
				8'h33 : r_dout <= #DLY 32'h4981ac83;
				8'h34 : r_dout <= #DLY 32'h334266ce;
				8'h35 : r_dout <= #DLY 32'h8c9341b7;
				8'h36 : r_dout <= #DLY 32'hd0d854c0;
				8'h37 : r_dout <= #DLY 32'hcb3a6c88;
				8'h38 : r_dout <= #DLY 32'h47bc2829;
				8'h39 : r_dout <= #DLY 32'h4725ba37;
				8'h3a : r_dout <= #DLY 32'ha66ad22b;
				8'h3b : r_dout <= #DLY 32'h7ad61f1e;
				8'h3c : r_dout <= #DLY 32'h0c5cbafa;
				8'h3d : r_dout <= #DLY 32'h4437f107;
				8'h3e : r_dout <= #DLY 32'hb6e79962;
				8'h3f : r_dout <= #DLY 32'h42d2d816;
				8'h40 : r_dout <= #DLY 32'h0a961288;
				8'h41 : r_dout <= #DLY 32'he1a5c06e;
				8'h42 : r_dout <= #DLY 32'h13749e67;
				8'h43 : r_dout <= #DLY 32'h72fc081a;
				8'h44 : r_dout <= #DLY 32'hb1d139f7;
				8'h45 : r_dout <= #DLY 32'hf9583745;
				8'h46 : r_dout <= #DLY 32'hcf19df58;
				8'h47 : r_dout <= #DLY 32'hbec3f756;
				8'h48 : r_dout <= #DLY 32'hc06eba30;
				8'h49 : r_dout <= #DLY 32'h07211b24;
				8'h4a : r_dout <= #DLY 32'h45c28829;
				8'h4b : r_dout <= #DLY 32'hc95e317f;
				8'h4c : r_dout <= #DLY 32'hbc8ec511;
				8'h4d : r_dout <= #DLY 32'h38bc46e9;
				8'h4e : r_dout <= #DLY 32'hc6e6fa14;
				8'h4f : r_dout <= #DLY 32'hbae8584a;
				8'h50 : r_dout <= #DLY 32'had4ebc46;
				8'h51 : r_dout <= #DLY 32'h468f508b;
				8'h52 : r_dout <= #DLY 32'h7829435f;
				8'h53 : r_dout <= #DLY 32'hf124183b;
				8'h54 : r_dout <= #DLY 32'h821dba9f;
				8'h55 : r_dout <= #DLY 32'haff60ff4;
				8'h56 : r_dout <= #DLY 32'hea2c4e6d;
				8'h57 : r_dout <= #DLY 32'h16e39264;
				8'h58 : r_dout <= #DLY 32'h92544a8b;
				8'h59 : r_dout <= #DLY 32'h009b4fc3;
				8'h5a : r_dout <= #DLY 32'haba68ced;
				8'h5b : r_dout <= #DLY 32'h9ac96f78;
				8'h5c : r_dout <= #DLY 32'h06a5b79a;
				8'h5d : r_dout <= #DLY 32'hb2856e6e;
				8'h5e : r_dout <= #DLY 32'h1aec3ca9;
				8'h5f : r_dout <= #DLY 32'hbe838688;
				8'h60 : r_dout <= #DLY 32'h0e0804e9;
				8'h61 : r_dout <= #DLY 32'h55f1be56;
				8'h62 : r_dout <= #DLY 32'he7e5363b;
				8'h63 : r_dout <= #DLY 32'hb3a1f25d;
				8'h64 : r_dout <= #DLY 32'hf7debb85;
				8'h65 : r_dout <= #DLY 32'h61fe033c;
				8'h66 : r_dout <= #DLY 32'h16746233;
				8'h67 : r_dout <= #DLY 32'h3c034c28;
				8'h68 : r_dout <= #DLY 32'hda6d0c74;
				8'h69 : r_dout <= #DLY 32'h79aac56c;
				8'h6a : r_dout <= #DLY 32'h3ce4e1ad;
				8'h6b : r_dout <= #DLY 32'h51f0c802;
				8'h6c : r_dout <= #DLY 32'h98f8f35a;
				8'h6d : r_dout <= #DLY 32'h1626a49f;
				8'h6e : r_dout <= #DLY 32'heed82b29;
				8'h6f : r_dout <= #DLY 32'h1d382fe3;
				8'h70 : r_dout <= #DLY 32'h0c4fb99a;
				8'h71 : r_dout <= #DLY 32'hbb325778;
				8'h72 : r_dout <= #DLY 32'h3ec6d97b;
				8'h73 : r_dout <= #DLY 32'h6e77a6a9;
				8'h74 : r_dout <= #DLY 32'hcb658b5c;
				8'h75 : r_dout <= #DLY 32'hd45230c7;
				8'h76 : r_dout <= #DLY 32'h2bd1408b;
				8'h77 : r_dout <= #DLY 32'h60c03eb7;
				8'h78 : r_dout <= #DLY 32'hb9068d78;
				8'h79 : r_dout <= #DLY 32'ha33754f4;
				8'h7a : r_dout <= #DLY 32'hf430c87d;
				8'h7b : r_dout <= #DLY 32'hc8a71302;
				8'h7c : r_dout <= #DLY 32'hb96d8c32;
				8'h7d : r_dout <= #DLY 32'hebd4e7be;
				8'h7e : r_dout <= #DLY 32'hbe8b9d2d;
				8'h7f : r_dout <= #DLY 32'h7979fb06;
				8'h80 : r_dout <= #DLY 32'he7225308;
				8'h81 : r_dout <= #DLY 32'h8b75cf77;
				8'h82 : r_dout <= #DLY 32'h11ef8da4;
				8'h83 : r_dout <= #DLY 32'he083c858;
				8'h84 : r_dout <= #DLY 32'h8d6b786f;
				8'h85 : r_dout <= #DLY 32'h5a6317a6;
				8'h86 : r_dout <= #DLY 32'hfa5cf7a0;
				8'h87 : r_dout <= #DLY 32'h5dda0033;
				8'h88 : r_dout <= #DLY 32'hf28ebfb0;
				8'h89 : r_dout <= #DLY 32'hf5b9c310;
				8'h8a : r_dout <= #DLY 32'ha0eac280;
				8'h8b : r_dout <= #DLY 32'h08b9767a;
				8'h8c : r_dout <= #DLY 32'ha3d9d2b0;
				8'h8d : r_dout <= #DLY 32'h79d34217;
				8'h8e : r_dout <= #DLY 32'h021a718d;
				8'h8f : r_dout <= #DLY 32'h9ac6336a;
				8'h90 : r_dout <= #DLY 32'h2711fd60;
				8'h91 : r_dout <= #DLY 32'h438050e3;
				8'h92 : r_dout <= #DLY 32'h069908a8;
				8'h93 : r_dout <= #DLY 32'h3d7fedc4;
				8'h94 : r_dout <= #DLY 32'h826d2bef;
				8'h95 : r_dout <= #DLY 32'h4eeb8476;
				8'h96 : r_dout <= #DLY 32'h488dcf25;
				8'h97 : r_dout <= #DLY 32'h36c9d566;
				8'h98 : r_dout <= #DLY 32'h28e74e41;
				8'h99 : r_dout <= #DLY 32'hc2610aca;
				8'h9a : r_dout <= #DLY 32'h3d49a9cf;
				8'h9b : r_dout <= #DLY 32'hbae3b9df;
				8'h9c : r_dout <= #DLY 32'hb65f8de6;
				8'h9d : r_dout <= #DLY 32'h92aeaf64;
				8'h9e : r_dout <= #DLY 32'h3ac7d5e6;
				8'h9f : r_dout <= #DLY 32'h9ea80509;
				8'ha0 : r_dout <= #DLY 32'hf22b017d;
				8'ha1 : r_dout <= #DLY 32'ha4173f70;
				8'ha2 : r_dout <= #DLY 32'hdd1e16c3;
				8'ha3 : r_dout <= #DLY 32'h15e0d7f9;
				8'ha4 : r_dout <= #DLY 32'h50b1b887;
				8'ha5 : r_dout <= #DLY 32'h2b9f4fd5;
				8'ha6 : r_dout <= #DLY 32'h625aba82;
				8'ha7 : r_dout <= #DLY 32'h6a017962;
				8'ha8 : r_dout <= #DLY 32'h2ec01b9c;
				8'ha9 : r_dout <= #DLY 32'h15488aa9;
				8'haa : r_dout <= #DLY 32'hd716e740;
				8'hab : r_dout <= #DLY 32'h40055a2c;
				8'hac : r_dout <= #DLY 32'h93d29a22;
				8'had : r_dout <= #DLY 32'he32dbf9a;
				8'hae : r_dout <= #DLY 32'h058745b9;
				8'haf : r_dout <= #DLY 32'h3453dc1e;
				8'hb0 : r_dout <= #DLY 32'hd699296e;
				8'hb1 : r_dout <= #DLY 32'h496cff6f;
				8'hb2 : r_dout <= #DLY 32'h1c9f4986;
				8'hb3 : r_dout <= #DLY 32'hdfe2ed07;
				8'hb4 : r_dout <= #DLY 32'hb87242d1;
				8'hb5 : r_dout <= #DLY 32'h19de7eae;
				8'hb6 : r_dout <= #DLY 32'h053e561a;
				8'hb7 : r_dout <= #DLY 32'h15ad6f8c;
				8'hb8 : r_dout <= #DLY 32'h66626c1c;
				8'hb9 : r_dout <= #DLY 32'h7154c24c;
				8'hba : r_dout <= #DLY 32'hea082b2a;
				8'hbb : r_dout <= #DLY 32'h93eb2939;
				8'hbc : r_dout <= #DLY 32'h17dcb0f0;
				8'hbd : r_dout <= #DLY 32'h58d4f2ae;
				8'hbe : r_dout <= #DLY 32'h9ea294fb;
				8'hbf : r_dout <= #DLY 32'h52cf564c;
				8'hc0 : r_dout <= #DLY 32'h9883fe66;
				8'hc1 : r_dout <= #DLY 32'h2ec40581;
				8'hc2 : r_dout <= #DLY 32'h763953c3;
				8'hc3 : r_dout <= #DLY 32'h01d6692e;
				8'hc4 : r_dout <= #DLY 32'hd3a0c108;
				8'hc5 : r_dout <= #DLY 32'ha1e7160e;
				8'hc6 : r_dout <= #DLY 32'he4f2dfa6;
				8'hc7 : r_dout <= #DLY 32'h693ed285;
				8'hc8 : r_dout <= #DLY 32'h74904698;
				8'hc9 : r_dout <= #DLY 32'h4c2b0edd;
				8'hca : r_dout <= #DLY 32'h4f757656;
				8'hcb : r_dout <= #DLY 32'h5d393378;
				8'hcc : r_dout <= #DLY 32'ha132234f;
				8'hcd : r_dout <= #DLY 32'h3d321c5d;
				8'hce : r_dout <= #DLY 32'hc3f5e194;
				8'hcf : r_dout <= #DLY 32'h4b269301;
				8'hd0 : r_dout <= #DLY 32'hc79f022f;
				8'hd1 : r_dout <= #DLY 32'h3c997e7e;
				8'hd2 : r_dout <= #DLY 32'h5e4f9504;
				8'hd3 : r_dout <= #DLY 32'h3ffafbbd;
				8'hd4 : r_dout <= #DLY 32'h76f7ad0e;
				8'hd5 : r_dout <= #DLY 32'h296693f4;
				8'hd6 : r_dout <= #DLY 32'h3d1fce6f;
				8'hd7 : r_dout <= #DLY 32'hc61e45be;
				8'hd8 : r_dout <= #DLY 32'hd3b5ab34;
				8'hd9 : r_dout <= #DLY 32'hf72bf9b7;
				8'hda : r_dout <= #DLY 32'h1b0434c0;
				8'hdb : r_dout <= #DLY 32'h4e72b567;
				8'hdc : r_dout <= #DLY 32'h5592a33d;
				8'hdd : r_dout <= #DLY 32'hb5229301;
				8'hde : r_dout <= #DLY 32'hcfd2a87f;
				8'hdf : r_dout <= #DLY 32'h60aeb767;
				8'he0 : r_dout <= #DLY 32'h1814386b;
				8'he1 : r_dout <= #DLY 32'h30bcc33d;
				8'he2 : r_dout <= #DLY 32'h38a0c07d;
				8'he3 : r_dout <= #DLY 32'hfd1606f2;
				8'he4 : r_dout <= #DLY 32'hc363519b;
				8'he5 : r_dout <= #DLY 32'h589dd390;
				8'he6 : r_dout <= #DLY 32'h5479f8e6;
				8'he7 : r_dout <= #DLY 32'h1cb8d647;
				8'he8 : r_dout <= #DLY 32'h97fd61a9;
				8'he9 : r_dout <= #DLY 32'hea7759f4;
				8'hea : r_dout <= #DLY 32'h2d57539d;
				8'heb : r_dout <= #DLY 32'h569a58cf;
				8'hec : r_dout <= #DLY 32'he84e63ad;
				8'hed : r_dout <= #DLY 32'h462e1b78;
				8'hee : r_dout <= #DLY 32'h6580f87e;
				8'hef : r_dout <= #DLY 32'hf3817914;
				8'hf0 : r_dout <= #DLY 32'h91da55f4;
				8'hf1 : r_dout <= #DLY 32'h40a230f3;
				8'hf2 : r_dout <= #DLY 32'hd1988f35;
				8'hf3 : r_dout <= #DLY 32'hb6e318d2;
				8'hf4 : r_dout <= #DLY 32'h3ffa50bc;
				8'hf5 : r_dout <= #DLY 32'h3d40f021;
				8'hf6 : r_dout <= #DLY 32'hc3c0bdae;
				8'hf7 : r_dout <= #DLY 32'h4958c24c;
				8'hf8 : r_dout <= #DLY 32'h518f36b2;
				8'hf9 : r_dout <= #DLY 32'h84b1d370;
				8'hfa : r_dout <= #DLY 32'h0fedce83;
				8'hfb : r_dout <= #DLY 32'h878ddada;
				8'hfc : r_dout <= #DLY 32'hf2a279c7;
				8'hfd : r_dout <= #DLY 32'h94e01be8;
				8'hfe : r_dout <= #DLY 32'h90716f4b;
				8'hff : r_dout <= #DLY 32'h954b8aa3;
			endcase
		end
    end

endmodule
