/*  
Copyright 2019 XCrypt Studio                
																	 
Licensed under the Apache License, Version 2.0 (the "License");         
you may not use this file except in compliance with the License.        
You may obtain a copy of the License at                                 
																	 
 http://www.apache.org/licenses/LICENSE-2.0                          
																	 
Unless required by applicable law or agreed to in writing, software    
distributed under the License is distributed on an "AS IS" BASIS,       
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and     
limitations under the License.                                          
*/  

// ------------------------------------------------------------------------------
// File name        :   cast5_sbox26.v
// Function         :   CAST5 Cryptographic Algorithm Core SBox-2 & SBox-6
// ------------------------------------------------------------------------------
// Author           :   Xie
// Version          ：  v-1.0
// Date				:   2019-2-2
// Email            :   xcrypt@126.com
// ------------------------------------------------------------------------------

`timescale 1ns / 1ps

module cast5_sbox26(
	input 			i_clk,
	input 			i_sel, //1: s-box 2 0:s-box 6
    input   [7:0]   i_addr,
    output  [31:0]  o_data
    );
	
	localparam DLY = 1;
	
    reg [31:0] r_dout;
    assign o_data = r_dout;
	//
    always@(posedge i_clk) begin
		if(i_sel) begin  
			case(i_addr)	//s-box 2
				8'h00 : r_dout <= #DLY 32'h1f201094;
				8'h01 : r_dout <= #DLY 32'hef0ba75b;
				8'h02 : r_dout <= #DLY 32'h69e3cf7e;
				8'h03 : r_dout <= #DLY 32'h393f4380;
				8'h04 : r_dout <= #DLY 32'hfe61cf7a;
				8'h05 : r_dout <= #DLY 32'heec5207a;
				8'h06 : r_dout <= #DLY 32'h55889c94;
				8'h07 : r_dout <= #DLY 32'h72fc0651;
				8'h08 : r_dout <= #DLY 32'hada7ef79;
				8'h09 : r_dout <= #DLY 32'h4e1d7235;
				8'h0a : r_dout <= #DLY 32'hd55a63ce;
				8'h0b : r_dout <= #DLY 32'hde0436ba;
				8'h0c : r_dout <= #DLY 32'h99c430ef;
				8'h0d : r_dout <= #DLY 32'h5f0c0794;
				8'h0e : r_dout <= #DLY 32'h18dcdb7d;
				8'h0f : r_dout <= #DLY 32'ha1d6eff3;
				8'h10 : r_dout <= #DLY 32'ha0b52f7b;
				8'h11 : r_dout <= #DLY 32'h59e83605;
				8'h12 : r_dout <= #DLY 32'hee15b094;
				8'h13 : r_dout <= #DLY 32'he9ffd909;
				8'h14 : r_dout <= #DLY 32'hdc440086;
				8'h15 : r_dout <= #DLY 32'hef944459;
				8'h16 : r_dout <= #DLY 32'hba83ccb3;
				8'h17 : r_dout <= #DLY 32'he0c3cdfb;
				8'h18 : r_dout <= #DLY 32'hd1da4181;
				8'h19 : r_dout <= #DLY 32'h3b092ab1;
				8'h1a : r_dout <= #DLY 32'hf997f1c1;
				8'h1b : r_dout <= #DLY 32'ha5e6cf7b;
				8'h1c : r_dout <= #DLY 32'h01420ddb;
				8'h1d : r_dout <= #DLY 32'he4e7ef5b;
				8'h1e : r_dout <= #DLY 32'h25a1ff41;
				8'h1f : r_dout <= #DLY 32'he180f806;
				8'h20 : r_dout <= #DLY 32'h1fc41080;
				8'h21 : r_dout <= #DLY 32'h179bee7a;
				8'h22 : r_dout <= #DLY 32'hd37ac6a9;
				8'h23 : r_dout <= #DLY 32'hfe5830a4;
				8'h24 : r_dout <= #DLY 32'h98de8b7f;
				8'h25 : r_dout <= #DLY 32'h77e83f4e;
				8'h26 : r_dout <= #DLY 32'h79929269;
				8'h27 : r_dout <= #DLY 32'h24fa9f7b;
				8'h28 : r_dout <= #DLY 32'he113c85b;
				8'h29 : r_dout <= #DLY 32'hacc40083;
				8'h2a : r_dout <= #DLY 32'hd7503525;
				8'h2b : r_dout <= #DLY 32'hf7ea615f;
				8'h2c : r_dout <= #DLY 32'h62143154;
				8'h2d : r_dout <= #DLY 32'h0d554b63;
				8'h2e : r_dout <= #DLY 32'h5d681121;
				8'h2f : r_dout <= #DLY 32'hc866c359;
				8'h30 : r_dout <= #DLY 32'h3d63cf73;
				8'h31 : r_dout <= #DLY 32'hcee234c0;
				8'h32 : r_dout <= #DLY 32'hd4d87e87;
				8'h33 : r_dout <= #DLY 32'h5c672b21;
				8'h34 : r_dout <= #DLY 32'h071f6181;
				8'h35 : r_dout <= #DLY 32'h39f7627f;
				8'h36 : r_dout <= #DLY 32'h361e3084;
				8'h37 : r_dout <= #DLY 32'he4eb573b;
				8'h38 : r_dout <= #DLY 32'h602f64a4;
				8'h39 : r_dout <= #DLY 32'hd63acd9c;
				8'h3a : r_dout <= #DLY 32'h1bbc4635;
				8'h3b : r_dout <= #DLY 32'h9e81032d;
				8'h3c : r_dout <= #DLY 32'h2701f50c;
				8'h3d : r_dout <= #DLY 32'h99847ab4;
				8'h3e : r_dout <= #DLY 32'ha0e3df79;
				8'h3f : r_dout <= #DLY 32'hba6cf38c;
				8'h40 : r_dout <= #DLY 32'h10843094;
				8'h41 : r_dout <= #DLY 32'h2537a95e;
				8'h42 : r_dout <= #DLY 32'hf46f6ffe;
				8'h43 : r_dout <= #DLY 32'ha1ff3b1f;
				8'h44 : r_dout <= #DLY 32'h208cfb6a;
				8'h45 : r_dout <= #DLY 32'h8f458c74;
				8'h46 : r_dout <= #DLY 32'hd9e0a227;
				8'h47 : r_dout <= #DLY 32'h4ec73a34;
				8'h48 : r_dout <= #DLY 32'hfc884f69;
				8'h49 : r_dout <= #DLY 32'h3e4de8df;
				8'h4a : r_dout <= #DLY 32'hef0e0088;
				8'h4b : r_dout <= #DLY 32'h3559648d;
				8'h4c : r_dout <= #DLY 32'h8a45388c;
				8'h4d : r_dout <= #DLY 32'h1d804366;
				8'h4e : r_dout <= #DLY 32'h721d9bfd;
				8'h4f : r_dout <= #DLY 32'ha58684bb;
				8'h50 : r_dout <= #DLY 32'he8256333;
				8'h51 : r_dout <= #DLY 32'h844e8212;
				8'h52 : r_dout <= #DLY 32'h128d8098;
				8'h53 : r_dout <= #DLY 32'hfed33fb4;
				8'h54 : r_dout <= #DLY 32'hce280ae1;
				8'h55 : r_dout <= #DLY 32'h27e19ba5;
				8'h56 : r_dout <= #DLY 32'hd5a6c252;
				8'h57 : r_dout <= #DLY 32'he49754bd;
				8'h58 : r_dout <= #DLY 32'hc5d655dd;
				8'h59 : r_dout <= #DLY 32'heb667064;
				8'h5a : r_dout <= #DLY 32'h77840b4d;
				8'h5b : r_dout <= #DLY 32'ha1b6a801;
				8'h5c : r_dout <= #DLY 32'h84db26a9;
				8'h5d : r_dout <= #DLY 32'he0b56714;
				8'h5e : r_dout <= #DLY 32'h21f043b7;
				8'h5f : r_dout <= #DLY 32'he5d05860;
				8'h60 : r_dout <= #DLY 32'h54f03084;
				8'h61 : r_dout <= #DLY 32'h066ff472;
				8'h62 : r_dout <= #DLY 32'ha31aa153;
				8'h63 : r_dout <= #DLY 32'hdadc4755;
				8'h64 : r_dout <= #DLY 32'hb5625dbf;
				8'h65 : r_dout <= #DLY 32'h68561be6;
				8'h66 : r_dout <= #DLY 32'h83ca6b94;
				8'h67 : r_dout <= #DLY 32'h2d6ed23b;
				8'h68 : r_dout <= #DLY 32'heccf01db;
				8'h69 : r_dout <= #DLY 32'ha6d3d0ba;
				8'h6a : r_dout <= #DLY 32'hb6803d5c;
				8'h6b : r_dout <= #DLY 32'haf77a709;
				8'h6c : r_dout <= #DLY 32'h33b4a34c;
				8'h6d : r_dout <= #DLY 32'h397bc8d6;
				8'h6e : r_dout <= #DLY 32'h5ee22b95;
				8'h6f : r_dout <= #DLY 32'h5f0e5304;
				8'h70 : r_dout <= #DLY 32'h81ed6f61;
				8'h71 : r_dout <= #DLY 32'h20e74364;
				8'h72 : r_dout <= #DLY 32'hb45e1378;
				8'h73 : r_dout <= #DLY 32'hde18639b;
				8'h74 : r_dout <= #DLY 32'h881ca122;
				8'h75 : r_dout <= #DLY 32'hb96726d1;
				8'h76 : r_dout <= #DLY 32'h8049a7e8;
				8'h77 : r_dout <= #DLY 32'h22b7da7b;
				8'h78 : r_dout <= #DLY 32'h5e552d25;
				8'h79 : r_dout <= #DLY 32'h5272d237;
				8'h7a : r_dout <= #DLY 32'h79d2951c;
				8'h7b : r_dout <= #DLY 32'hc60d894c;
				8'h7c : r_dout <= #DLY 32'h488cb402;
				8'h7d : r_dout <= #DLY 32'h1ba4fe5b;
				8'h7e : r_dout <= #DLY 32'ha4b09f6b;
				8'h7f : r_dout <= #DLY 32'h1ca815cf;
				8'h80 : r_dout <= #DLY 32'ha20c3005;
				8'h81 : r_dout <= #DLY 32'h8871df63;
				8'h82 : r_dout <= #DLY 32'hb9de2fcb;
				8'h83 : r_dout <= #DLY 32'h0cc6c9e9;
				8'h84 : r_dout <= #DLY 32'h0beeff53;
				8'h85 : r_dout <= #DLY 32'he3214517;
				8'h86 : r_dout <= #DLY 32'hb4542835;
				8'h87 : r_dout <= #DLY 32'h9f63293c;
				8'h88 : r_dout <= #DLY 32'hee41e729;
				8'h89 : r_dout <= #DLY 32'h6e1d2d7c;
				8'h8a : r_dout <= #DLY 32'h50045286;
				8'h8b : r_dout <= #DLY 32'h1e6685f3;
				8'h8c : r_dout <= #DLY 32'hf33401c6;
				8'h8d : r_dout <= #DLY 32'h30a22c95;
				8'h8e : r_dout <= #DLY 32'h31a70850;
				8'h8f : r_dout <= #DLY 32'h60930f13;
				8'h90 : r_dout <= #DLY 32'h73f98417;
				8'h91 : r_dout <= #DLY 32'ha1269859;
				8'h92 : r_dout <= #DLY 32'hec645c44;
				8'h93 : r_dout <= #DLY 32'h52c877a9;
				8'h94 : r_dout <= #DLY 32'hcdff33a6;
				8'h95 : r_dout <= #DLY 32'ha02b1741;
				8'h96 : r_dout <= #DLY 32'h7cbad9a2;
				8'h97 : r_dout <= #DLY 32'h2180036f;
				8'h98 : r_dout <= #DLY 32'h50d99c08;
				8'h99 : r_dout <= #DLY 32'hcb3f4861;
				8'h9a : r_dout <= #DLY 32'hc26bd765;
				8'h9b : r_dout <= #DLY 32'h64a3f6ab;
				8'h9c : r_dout <= #DLY 32'h80342676;
				8'h9d : r_dout <= #DLY 32'h25a75e7b;
				8'h9e : r_dout <= #DLY 32'he4e6d1fc;
				8'h9f : r_dout <= #DLY 32'h20c710e6;
				8'ha0 : r_dout <= #DLY 32'hcdf0b680;
				8'ha1 : r_dout <= #DLY 32'h17844d3b;
				8'ha2 : r_dout <= #DLY 32'h31eef84d;
				8'ha3 : r_dout <= #DLY 32'h7e0824e4;
				8'ha4 : r_dout <= #DLY 32'h2ccb49eb;
				8'ha5 : r_dout <= #DLY 32'h846a3bae;
				8'ha6 : r_dout <= #DLY 32'h8ff77888;
				8'ha7 : r_dout <= #DLY 32'hee5d60f6;
				8'ha8 : r_dout <= #DLY 32'h7af75673;
				8'ha9 : r_dout <= #DLY 32'h2fdd5cdb;
				8'haa : r_dout <= #DLY 32'ha11631c1;
				8'hab : r_dout <= #DLY 32'h30f66f43;
				8'hac : r_dout <= #DLY 32'hb3faec54;
				8'had : r_dout <= #DLY 32'h157fd7fa;
				8'hae : r_dout <= #DLY 32'hef8579cc;
				8'haf : r_dout <= #DLY 32'hd152de58;
				8'hb0 : r_dout <= #DLY 32'hdb2ffd5e;
				8'hb1 : r_dout <= #DLY 32'h8f32ce19;
				8'hb2 : r_dout <= #DLY 32'h306af97a;
				8'hb3 : r_dout <= #DLY 32'h02f03ef8;
				8'hb4 : r_dout <= #DLY 32'h99319ad5;
				8'hb5 : r_dout <= #DLY 32'hc242fa0f;
				8'hb6 : r_dout <= #DLY 32'ha7e3ebb0;
				8'hb7 : r_dout <= #DLY 32'hc68e4906;
				8'hb8 : r_dout <= #DLY 32'hb8da230c;
				8'hb9 : r_dout <= #DLY 32'h80823028;
				8'hba : r_dout <= #DLY 32'hdcdef3c8;
				8'hbb : r_dout <= #DLY 32'hd35fb171;
				8'hbc : r_dout <= #DLY 32'h088a1bc8;
				8'hbd : r_dout <= #DLY 32'hbec0c560;
				8'hbe : r_dout <= #DLY 32'h61a3c9e8;
				8'hbf : r_dout <= #DLY 32'hbca8f54d;
				8'hc0 : r_dout <= #DLY 32'hc72feffa;
				8'hc1 : r_dout <= #DLY 32'h22822e99;
				8'hc2 : r_dout <= #DLY 32'h82c570b4;
				8'hc3 : r_dout <= #DLY 32'hd8d94e89;
				8'hc4 : r_dout <= #DLY 32'h8b1c34bc;
				8'hc5 : r_dout <= #DLY 32'h301e16e6;
				8'hc6 : r_dout <= #DLY 32'h273be979;
				8'hc7 : r_dout <= #DLY 32'hb0ffeaa6;
				8'hc8 : r_dout <= #DLY 32'h61d9b8c6;
				8'hc9 : r_dout <= #DLY 32'h00b24869;
				8'hca : r_dout <= #DLY 32'hb7ffce3f;
				8'hcb : r_dout <= #DLY 32'h08dc283b;
				8'hcc : r_dout <= #DLY 32'h43daf65a;
				8'hcd : r_dout <= #DLY 32'hf7e19798;
				8'hce : r_dout <= #DLY 32'h7619b72f;
				8'hcf : r_dout <= #DLY 32'h8f1c9ba4;
				8'hd0 : r_dout <= #DLY 32'hdc8637a0;
				8'hd1 : r_dout <= #DLY 32'h16a7d3b1;
				8'hd2 : r_dout <= #DLY 32'h9fc393b7;
				8'hd3 : r_dout <= #DLY 32'ha7136eeb;
				8'hd4 : r_dout <= #DLY 32'hc6bcc63e;
				8'hd5 : r_dout <= #DLY 32'h1a513742;
				8'hd6 : r_dout <= #DLY 32'hef6828bc;
				8'hd7 : r_dout <= #DLY 32'h520365d6;
				8'hd8 : r_dout <= #DLY 32'h2d6a77ab;
				8'hd9 : r_dout <= #DLY 32'h3527ed4b;
				8'hda : r_dout <= #DLY 32'h821fd216;
				8'hdb : r_dout <= #DLY 32'h095c6e2e;
				8'hdc : r_dout <= #DLY 32'hdb92f2fb;
				8'hdd : r_dout <= #DLY 32'h5eea29cb;
				8'hde : r_dout <= #DLY 32'h145892f5;
				8'hdf : r_dout <= #DLY 32'h91584f7f;
				8'he0 : r_dout <= #DLY 32'h5483697b;
				8'he1 : r_dout <= #DLY 32'h2667a8cc;
				8'he2 : r_dout <= #DLY 32'h85196048;
				8'he3 : r_dout <= #DLY 32'h8c4bacea;
				8'he4 : r_dout <= #DLY 32'h833860d4;
				8'he5 : r_dout <= #DLY 32'h0d23e0f9;
				8'he6 : r_dout <= #DLY 32'h6c387e8a;
				8'he7 : r_dout <= #DLY 32'h0ae6d249;
				8'he8 : r_dout <= #DLY 32'hb284600c;
				8'he9 : r_dout <= #DLY 32'hd835731d;
				8'hea : r_dout <= #DLY 32'hdcb1c647;
				8'heb : r_dout <= #DLY 32'hac4c56ea;
				8'hec : r_dout <= #DLY 32'h3ebd81b3;
				8'hed : r_dout <= #DLY 32'h230eabb0;
				8'hee : r_dout <= #DLY 32'h6438bc87;
				8'hef : r_dout <= #DLY 32'hf0b5b1fa;
				8'hf0 : r_dout <= #DLY 32'h8f5ea2b3;
				8'hf1 : r_dout <= #DLY 32'hfc184642;
				8'hf2 : r_dout <= #DLY 32'h0a036b7a;
				8'hf3 : r_dout <= #DLY 32'h4fb089bd;
				8'hf4 : r_dout <= #DLY 32'h649da589;
				8'hf5 : r_dout <= #DLY 32'ha345415e;
				8'hf6 : r_dout <= #DLY 32'h5c038323;
				8'hf7 : r_dout <= #DLY 32'h3e5d3bb9;
				8'hf8 : r_dout <= #DLY 32'h43d79572;
				8'hf9 : r_dout <= #DLY 32'h7e6dd07c;
				8'hfa : r_dout <= #DLY 32'h06dfdf1e;
				8'hfb : r_dout <= #DLY 32'h6c6cc4ef;
				8'hfc : r_dout <= #DLY 32'h7160a539;
				8'hfd : r_dout <= #DLY 32'h73bfbe70;
				8'hfe : r_dout <= #DLY 32'h83877605;
				8'hff : r_dout <= #DLY 32'h4523ecf1;
			endcase
		end else begin    
			case(i_addr)	//s-box 6
				8'h00 : r_dout <= #DLY 32'hf6fa8f9d;
				8'h01 : r_dout <= #DLY 32'h2cac6ce1;
				8'h02 : r_dout <= #DLY 32'h4ca34867;
				8'h03 : r_dout <= #DLY 32'he2337f7c;
				8'h04 : r_dout <= #DLY 32'h95db08e7;
				8'h05 : r_dout <= #DLY 32'h016843b4;
				8'h06 : r_dout <= #DLY 32'heced5cbc;
				8'h07 : r_dout <= #DLY 32'h325553ac;
				8'h08 : r_dout <= #DLY 32'hbf9f0960;
				8'h09 : r_dout <= #DLY 32'hdfa1e2ed;
				8'h0a : r_dout <= #DLY 32'h83f0579d;
				8'h0b : r_dout <= #DLY 32'h63ed86b9;
				8'h0c : r_dout <= #DLY 32'h1ab6a6b8;
				8'h0d : r_dout <= #DLY 32'hde5ebe39;
				8'h0e : r_dout <= #DLY 32'hf38ff732;
				8'h0f : r_dout <= #DLY 32'h8989b138;
				8'h10 : r_dout <= #DLY 32'h33f14961;
				8'h11 : r_dout <= #DLY 32'hc01937bd;
				8'h12 : r_dout <= #DLY 32'hf506c6da;
				8'h13 : r_dout <= #DLY 32'he4625e7e;
				8'h14 : r_dout <= #DLY 32'ha308ea99;
				8'h15 : r_dout <= #DLY 32'h4e23e33c;
				8'h16 : r_dout <= #DLY 32'h79cbd7cc;
				8'h17 : r_dout <= #DLY 32'h48a14367;
				8'h18 : r_dout <= #DLY 32'ha3149619;
				8'h19 : r_dout <= #DLY 32'hfec94bd5;
				8'h1a : r_dout <= #DLY 32'ha114174a;
				8'h1b : r_dout <= #DLY 32'heaa01866;
				8'h1c : r_dout <= #DLY 32'ha084db2d;
				8'h1d : r_dout <= #DLY 32'h09a8486f;
				8'h1e : r_dout <= #DLY 32'ha888614a;
				8'h1f : r_dout <= #DLY 32'h2900af98;
				8'h20 : r_dout <= #DLY 32'h01665991;
				8'h21 : r_dout <= #DLY 32'he1992863;
				8'h22 : r_dout <= #DLY 32'hc8f30c60;
				8'h23 : r_dout <= #DLY 32'h2e78ef3c;
				8'h24 : r_dout <= #DLY 32'hd0d51932;
				8'h25 : r_dout <= #DLY 32'hcf0fec14;
				8'h26 : r_dout <= #DLY 32'hf7ca07d2;
				8'h27 : r_dout <= #DLY 32'hd0a82072;
				8'h28 : r_dout <= #DLY 32'hfd41197e;
				8'h29 : r_dout <= #DLY 32'h9305a6b0;
				8'h2a : r_dout <= #DLY 32'he86be3da;
				8'h2b : r_dout <= #DLY 32'h74bed3cd;
				8'h2c : r_dout <= #DLY 32'h372da53c;
				8'h2d : r_dout <= #DLY 32'h4c7f4448;
				8'h2e : r_dout <= #DLY 32'hdab5d440;
				8'h2f : r_dout <= #DLY 32'h6dba0ec3;
				8'h30 : r_dout <= #DLY 32'h083919a7;
				8'h31 : r_dout <= #DLY 32'h9fbaeed9;
				8'h32 : r_dout <= #DLY 32'h49dbcfb0;
				8'h33 : r_dout <= #DLY 32'h4e670c53;
				8'h34 : r_dout <= #DLY 32'h5c3d9c01;
				8'h35 : r_dout <= #DLY 32'h64bdb941;
				8'h36 : r_dout <= #DLY 32'h2c0e636a;
				8'h37 : r_dout <= #DLY 32'hba7dd9cd;
				8'h38 : r_dout <= #DLY 32'hea6f7388;
				8'h39 : r_dout <= #DLY 32'he70bc762;
				8'h3a : r_dout <= #DLY 32'h35f29adb;
				8'h3b : r_dout <= #DLY 32'h5c4cdd8d;
				8'h3c : r_dout <= #DLY 32'hf0d48d8c;
				8'h3d : r_dout <= #DLY 32'hb88153e2;
				8'h3e : r_dout <= #DLY 32'h08a19866;
				8'h3f : r_dout <= #DLY 32'h1ae2eac8;
				8'h40 : r_dout <= #DLY 32'h284caf89;
				8'h41 : r_dout <= #DLY 32'haa928223;
				8'h42 : r_dout <= #DLY 32'h9334be53;
				8'h43 : r_dout <= #DLY 32'h3b3a21bf;
				8'h44 : r_dout <= #DLY 32'h16434be3;
				8'h45 : r_dout <= #DLY 32'h9aea3906;
				8'h46 : r_dout <= #DLY 32'hefe8c36e;
				8'h47 : r_dout <= #DLY 32'hf890cdd9;
				8'h48 : r_dout <= #DLY 32'h80226dae;
				8'h49 : r_dout <= #DLY 32'hc340a4a3;
				8'h4a : r_dout <= #DLY 32'hdf7e9c09;
				8'h4b : r_dout <= #DLY 32'ha694a807;
				8'h4c : r_dout <= #DLY 32'h5b7c5ecc;
				8'h4d : r_dout <= #DLY 32'h221db3a6;
				8'h4e : r_dout <= #DLY 32'h9a69a02f;
				8'h4f : r_dout <= #DLY 32'h68818a54;
				8'h50 : r_dout <= #DLY 32'hceb2296f;
				8'h51 : r_dout <= #DLY 32'h53c0843a;
				8'h52 : r_dout <= #DLY 32'hfe893655;
				8'h53 : r_dout <= #DLY 32'h25bfe68a;
				8'h54 : r_dout <= #DLY 32'hb4628abc;
				8'h55 : r_dout <= #DLY 32'hcf222ebf;
				8'h56 : r_dout <= #DLY 32'h25ac6f48;
				8'h57 : r_dout <= #DLY 32'ha9a99387;
				8'h58 : r_dout <= #DLY 32'h53bddb65;
				8'h59 : r_dout <= #DLY 32'he76ffbe7;
				8'h5a : r_dout <= #DLY 32'he967fd78;
				8'h5b : r_dout <= #DLY 32'h0ba93563;
				8'h5c : r_dout <= #DLY 32'h8e342bc1;
				8'h5d : r_dout <= #DLY 32'he8a11be9;
				8'h5e : r_dout <= #DLY 32'h4980740d;
				8'h5f : r_dout <= #DLY 32'hc8087dfc;
				8'h60 : r_dout <= #DLY 32'h8de4bf99;
				8'h61 : r_dout <= #DLY 32'ha11101a0;
				8'h62 : r_dout <= #DLY 32'h7fd37975;
				8'h63 : r_dout <= #DLY 32'hda5a26c0;
				8'h64 : r_dout <= #DLY 32'he81f994f;
				8'h65 : r_dout <= #DLY 32'h9528cd89;
				8'h66 : r_dout <= #DLY 32'hfd339fed;
				8'h67 : r_dout <= #DLY 32'hb87834bf;
				8'h68 : r_dout <= #DLY 32'h5f04456d;
				8'h69 : r_dout <= #DLY 32'h22258698;
				8'h6a : r_dout <= #DLY 32'hc9c4c83b;
				8'h6b : r_dout <= #DLY 32'h2dc156be;
				8'h6c : r_dout <= #DLY 32'h4f628daa;
				8'h6d : r_dout <= #DLY 32'h57f55ec5;
				8'h6e : r_dout <= #DLY 32'he2220abe;
				8'h6f : r_dout <= #DLY 32'hd2916ebf;
				8'h70 : r_dout <= #DLY 32'h4ec75b95;
				8'h71 : r_dout <= #DLY 32'h24f2c3c0;
				8'h72 : r_dout <= #DLY 32'h42d15d99;
				8'h73 : r_dout <= #DLY 32'hcd0d7fa0;
				8'h74 : r_dout <= #DLY 32'h7b6e27ff;
				8'h75 : r_dout <= #DLY 32'ha8dc8af0;
				8'h76 : r_dout <= #DLY 32'h7345c106;
				8'h77 : r_dout <= #DLY 32'hf41e232f;
				8'h78 : r_dout <= #DLY 32'h35162386;
				8'h79 : r_dout <= #DLY 32'he6ea8926;
				8'h7a : r_dout <= #DLY 32'h3333b094;
				8'h7b : r_dout <= #DLY 32'h157ec6f2;
				8'h7c : r_dout <= #DLY 32'h372b74af;
				8'h7d : r_dout <= #DLY 32'h692573e4;
				8'h7e : r_dout <= #DLY 32'he9a9d848;
				8'h7f : r_dout <= #DLY 32'hf3160289;
				8'h80 : r_dout <= #DLY 32'h3a62ef1d;
				8'h81 : r_dout <= #DLY 32'ha787e238;
				8'h82 : r_dout <= #DLY 32'hf3a5f676;
				8'h83 : r_dout <= #DLY 32'h74364853;
				8'h84 : r_dout <= #DLY 32'h20951063;
				8'h85 : r_dout <= #DLY 32'h4576698d;
				8'h86 : r_dout <= #DLY 32'hb6fad407;
				8'h87 : r_dout <= #DLY 32'h592af950;
				8'h88 : r_dout <= #DLY 32'h36f73523;
				8'h89 : r_dout <= #DLY 32'h4cfb6e87;
				8'h8a : r_dout <= #DLY 32'h7da4cec0;
				8'h8b : r_dout <= #DLY 32'h6c152daa;
				8'h8c : r_dout <= #DLY 32'hcb0396a8;
				8'h8d : r_dout <= #DLY 32'hc50dfe5d;
				8'h8e : r_dout <= #DLY 32'hfcd707ab;
				8'h8f : r_dout <= #DLY 32'h0921c42f;
				8'h90 : r_dout <= #DLY 32'h89dff0bb;
				8'h91 : r_dout <= #DLY 32'h5fe2be78;
				8'h92 : r_dout <= #DLY 32'h448f4f33;
				8'h93 : r_dout <= #DLY 32'h754613c9;
				8'h94 : r_dout <= #DLY 32'h2b05d08d;
				8'h95 : r_dout <= #DLY 32'h48b9d585;
				8'h96 : r_dout <= #DLY 32'hdc049441;
				8'h97 : r_dout <= #DLY 32'hc8098f9b;
				8'h98 : r_dout <= #DLY 32'h7dede786;
				8'h99 : r_dout <= #DLY 32'hc39a3373;
				8'h9a : r_dout <= #DLY 32'h42410005;
				8'h9b : r_dout <= #DLY 32'h6a091751;
				8'h9c : r_dout <= #DLY 32'h0ef3c8a6;
				8'h9d : r_dout <= #DLY 32'h890072d6;
				8'h9e : r_dout <= #DLY 32'h28207682;
				8'h9f : r_dout <= #DLY 32'ha9a9f7be;
				8'ha0 : r_dout <= #DLY 32'hbf32679d;
				8'ha1 : r_dout <= #DLY 32'hd45b5b75;
				8'ha2 : r_dout <= #DLY 32'hb353fd00;
				8'ha3 : r_dout <= #DLY 32'hcbb0e358;
				8'ha4 : r_dout <= #DLY 32'h830f220a;
				8'ha5 : r_dout <= #DLY 32'h1f8fb214;
				8'ha6 : r_dout <= #DLY 32'hd372cf08;
				8'ha7 : r_dout <= #DLY 32'hcc3c4a13;
				8'ha8 : r_dout <= #DLY 32'h8cf63166;
				8'ha9 : r_dout <= #DLY 32'h061c87be;
				8'haa : r_dout <= #DLY 32'h88c98f88;
				8'hab : r_dout <= #DLY 32'h6062e397;
				8'hac : r_dout <= #DLY 32'h47cf8e7a;
				8'had : r_dout <= #DLY 32'hb6c85283;
				8'hae : r_dout <= #DLY 32'h3cc2acfb;
				8'haf : r_dout <= #DLY 32'h3fc06976;
				8'hb0 : r_dout <= #DLY 32'h4e8f0252;
				8'hb1 : r_dout <= #DLY 32'h64d8314d;
				8'hb2 : r_dout <= #DLY 32'hda3870e3;
				8'hb3 : r_dout <= #DLY 32'h1e665459;
				8'hb4 : r_dout <= #DLY 32'hc10908f0;
				8'hb5 : r_dout <= #DLY 32'h513021a5;
				8'hb6 : r_dout <= #DLY 32'h6c5b68b7;
				8'hb7 : r_dout <= #DLY 32'h822f8aa0;
				8'hb8 : r_dout <= #DLY 32'h3007cd3e;
				8'hb9 : r_dout <= #DLY 32'h74719eef;
				8'hba : r_dout <= #DLY 32'hdc872681;
				8'hbb : r_dout <= #DLY 32'h073340d4;
				8'hbc : r_dout <= #DLY 32'h7e432fd9;
				8'hbd : r_dout <= #DLY 32'h0c5ec241;
				8'hbe : r_dout <= #DLY 32'h8809286c;
				8'hbf : r_dout <= #DLY 32'hf592d891;
				8'hc0 : r_dout <= #DLY 32'h08a930f6;
				8'hc1 : r_dout <= #DLY 32'h957ef305;
				8'hc2 : r_dout <= #DLY 32'hb7fbffbd;
				8'hc3 : r_dout <= #DLY 32'hc266e96f;
				8'hc4 : r_dout <= #DLY 32'h6fe4ac98;
				8'hc5 : r_dout <= #DLY 32'hb173ecc0;
				8'hc6 : r_dout <= #DLY 32'hbc60b42a;
				8'hc7 : r_dout <= #DLY 32'h953498da;
				8'hc8 : r_dout <= #DLY 32'hfba1ae12;
				8'hc9 : r_dout <= #DLY 32'h2d4bd736;
				8'hca : r_dout <= #DLY 32'h0f25faab;
				8'hcb : r_dout <= #DLY 32'ha4f3fceb;
				8'hcc : r_dout <= #DLY 32'he2969123;
				8'hcd : r_dout <= #DLY 32'h257f0c3d;
				8'hce : r_dout <= #DLY 32'h9348af49;
				8'hcf : r_dout <= #DLY 32'h361400bc;
				8'hd0 : r_dout <= #DLY 32'he8816f4a;
				8'hd1 : r_dout <= #DLY 32'h3814f200;
				8'hd2 : r_dout <= #DLY 32'ha3f94043;
				8'hd3 : r_dout <= #DLY 32'h9c7a54c2;
				8'hd4 : r_dout <= #DLY 32'hbc704f57;
				8'hd5 : r_dout <= #DLY 32'hda41e7f9;
				8'hd6 : r_dout <= #DLY 32'hc25ad33a;
				8'hd7 : r_dout <= #DLY 32'h54f4a084;
				8'hd8 : r_dout <= #DLY 32'hb17f5505;
				8'hd9 : r_dout <= #DLY 32'h59357cbe;
				8'hda : r_dout <= #DLY 32'hedbd15c8;
				8'hdb : r_dout <= #DLY 32'h7f97c5ab;
				8'hdc : r_dout <= #DLY 32'hba5ac7b5;
				8'hdd : r_dout <= #DLY 32'hb6f6deaf;
				8'hde : r_dout <= #DLY 32'h3a479c3a;
				8'hdf : r_dout <= #DLY 32'h5302da25;
				8'he0 : r_dout <= #DLY 32'h653d7e6a;
				8'he1 : r_dout <= #DLY 32'h54268d49;
				8'he2 : r_dout <= #DLY 32'h51a477ea;
				8'he3 : r_dout <= #DLY 32'h5017d55b;
				8'he4 : r_dout <= #DLY 32'hd7d25d88;
				8'he5 : r_dout <= #DLY 32'h44136c76;
				8'he6 : r_dout <= #DLY 32'h0404a8c8;
				8'he7 : r_dout <= #DLY 32'hb8e5a121;
				8'he8 : r_dout <= #DLY 32'hb81a928a;
				8'he9 : r_dout <= #DLY 32'h60ed5869;
				8'hea : r_dout <= #DLY 32'h97c55b96;
				8'heb : r_dout <= #DLY 32'heaec991b;
				8'hec : r_dout <= #DLY 32'h29935913;
				8'hed : r_dout <= #DLY 32'h01fdb7f1;
				8'hee : r_dout <= #DLY 32'h088e8dfa;
				8'hef : r_dout <= #DLY 32'h9ab6f6f5;
				8'hf0 : r_dout <= #DLY 32'h3b4cbf9f;
				8'hf1 : r_dout <= #DLY 32'h4a5de3ab;
				8'hf2 : r_dout <= #DLY 32'he6051d35;
				8'hf3 : r_dout <= #DLY 32'ha0e1d855;
				8'hf4 : r_dout <= #DLY 32'hd36b4cf1;
				8'hf5 : r_dout <= #DLY 32'hf544edeb;
				8'hf6 : r_dout <= #DLY 32'hb0e93524;
				8'hf7 : r_dout <= #DLY 32'hbebb8fbd;
				8'hf8 : r_dout <= #DLY 32'ha2d762cf;
				8'hf9 : r_dout <= #DLY 32'h49c92f54;
				8'hfa : r_dout <= #DLY 32'h38b5f331;
				8'hfb : r_dout <= #DLY 32'h7128a454;
				8'hfc : r_dout <= #DLY 32'h48392905;
				8'hfd : r_dout <= #DLY 32'ha65b1db8;
				8'hfe : r_dout <= #DLY 32'h851c97bd;
				8'hff : r_dout <= #DLY 32'hd675cf2f;
			endcase
		end
	end

endmodule
