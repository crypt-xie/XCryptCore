/*  
Copyright 2019 XCrypt Studio                
																	 
Licensed under the Apache License, Version 2.0 (the "License");         
you may not use this file except in compliance with the License.        
You may obtain a copy of the License at                                 
																	 
 http://www.apache.org/licenses/LICENSE-2.0                          
																	 
Unless required by applicable law or agreed to in writing, software    
distributed under the License is distributed on an "AS IS" BASIS,       
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and     
limitations under the License.                                          
*/  

// ------------------------------------------------------------------------------
// File name        :   cast5_sbox4.v
// Function         :   CAST5 Cryptographic Algorithm Core SBox-4 & SBox-8
// ------------------------------------------------------------------------------
// Author           :   Xie
// Version          ：  v-1.0
// Date				:   2019-2-2
// Email            :   xcrypt@126.com
// ------------------------------------------------------------------------------

`timescale 1ns / 1ps

module cast5_sbox48(
	input 			i_clk,
	input			i_sel,  //1: s-box4 0:s-box8
    input   [7:0]   i_addr,
    output  [31:0]  o_data
    );
	
	localparam DLY = 1;
	
    reg [31:0] r_dout;
    assign o_data = r_dout;
	//
    always@(posedge i_clk) begin
		if(i_sel) begin  //s-box4
			case(i_addr)
				8'h00 : r_dout <= #DLY 32'h9db30420;
				8'h01 : r_dout <= #DLY 32'h1fb6e9de;
				8'h02 : r_dout <= #DLY 32'ha7be7bef;
				8'h03 : r_dout <= #DLY 32'hd273a298;
				8'h04 : r_dout <= #DLY 32'h4a4f7bdb;
				8'h05 : r_dout <= #DLY 32'h64ad8c57;
				8'h06 : r_dout <= #DLY 32'h85510443;
				8'h07 : r_dout <= #DLY 32'hfa020ed1;
				8'h08 : r_dout <= #DLY 32'h7e287aff;
				8'h09 : r_dout <= #DLY 32'he60fb663;
				8'h0a : r_dout <= #DLY 32'h095f35a1;
				8'h0b : r_dout <= #DLY 32'h79ebf120;
				8'h0c : r_dout <= #DLY 32'hfd059d43;
				8'h0d : r_dout <= #DLY 32'h6497b7b1;
				8'h0e : r_dout <= #DLY 32'hf3641f63;
				8'h0f : r_dout <= #DLY 32'h241e4adf;
				8'h10 : r_dout <= #DLY 32'h28147f5f;
				8'h11 : r_dout <= #DLY 32'h4fa2b8cd;
				8'h12 : r_dout <= #DLY 32'hc9430040;
				8'h13 : r_dout <= #DLY 32'h0cc32220;
				8'h14 : r_dout <= #DLY 32'hfdd30b30;
				8'h15 : r_dout <= #DLY 32'hc0a5374f;
				8'h16 : r_dout <= #DLY 32'h1d2d00d9;
				8'h17 : r_dout <= #DLY 32'h24147b15;
				8'h18 : r_dout <= #DLY 32'hee4d111a;
				8'h19 : r_dout <= #DLY 32'h0fca5167;
				8'h1a : r_dout <= #DLY 32'h71ff904c;
				8'h1b : r_dout <= #DLY 32'h2d195ffe;
				8'h1c : r_dout <= #DLY 32'h1a05645f;
				8'h1d : r_dout <= #DLY 32'h0c13fefe;
				8'h1e : r_dout <= #DLY 32'h081b08ca;
				8'h1f : r_dout <= #DLY 32'h05170121;
				8'h20 : r_dout <= #DLY 32'h80530100;
				8'h21 : r_dout <= #DLY 32'he83e5efe;
				8'h22 : r_dout <= #DLY 32'hac9af4f8;
				8'h23 : r_dout <= #DLY 32'h7fe72701;
				8'h24 : r_dout <= #DLY 32'hd2b8ee5f;
				8'h25 : r_dout <= #DLY 32'h06df4261;
				8'h26 : r_dout <= #DLY 32'hbb9e9b8a;
				8'h27 : r_dout <= #DLY 32'h7293ea25;
				8'h28 : r_dout <= #DLY 32'hce84ffdf;
				8'h29 : r_dout <= #DLY 32'hf5718801;
				8'h2a : r_dout <= #DLY 32'h3dd64b04;
				8'h2b : r_dout <= #DLY 32'ha26f263b;
				8'h2c : r_dout <= #DLY 32'h7ed48400;
				8'h2d : r_dout <= #DLY 32'h547eebe6;
				8'h2e : r_dout <= #DLY 32'h446d4ca0;
				8'h2f : r_dout <= #DLY 32'h6cf3d6f5;
				8'h30 : r_dout <= #DLY 32'h2649abdf;
				8'h31 : r_dout <= #DLY 32'haea0c7f5;
				8'h32 : r_dout <= #DLY 32'h36338cc1;
				8'h33 : r_dout <= #DLY 32'h503f7e93;
				8'h34 : r_dout <= #DLY 32'hd3772061;
				8'h35 : r_dout <= #DLY 32'h11b638e1;
				8'h36 : r_dout <= #DLY 32'h72500e03;
				8'h37 : r_dout <= #DLY 32'hf80eb2bb;
				8'h38 : r_dout <= #DLY 32'habe0502e;
				8'h39 : r_dout <= #DLY 32'hec8d77de;
				8'h3a : r_dout <= #DLY 32'h57971e81;
				8'h3b : r_dout <= #DLY 32'he14f6746;
				8'h3c : r_dout <= #DLY 32'hc9335400;
				8'h3d : r_dout <= #DLY 32'h6920318f;
				8'h3e : r_dout <= #DLY 32'h081dbb99;
				8'h3f : r_dout <= #DLY 32'hffc304a5;
				8'h40 : r_dout <= #DLY 32'h4d351805;
				8'h41 : r_dout <= #DLY 32'h7f3d5ce3;
				8'h42 : r_dout <= #DLY 32'ha6c866c6;
				8'h43 : r_dout <= #DLY 32'h5d5bcca9;
				8'h44 : r_dout <= #DLY 32'hdaec6fea;
				8'h45 : r_dout <= #DLY 32'h9f926f91;
				8'h46 : r_dout <= #DLY 32'h9f46222f;
				8'h47 : r_dout <= #DLY 32'h3991467d;
				8'h48 : r_dout <= #DLY 32'ha5bf6d8e;
				8'h49 : r_dout <= #DLY 32'h1143c44f;
				8'h4a : r_dout <= #DLY 32'h43958302;
				8'h4b : r_dout <= #DLY 32'hd0214eeb;
				8'h4c : r_dout <= #DLY 32'h022083b8;
				8'h4d : r_dout <= #DLY 32'h3fb6180c;
				8'h4e : r_dout <= #DLY 32'h18f8931e;
				8'h4f : r_dout <= #DLY 32'h281658e6;
				8'h50 : r_dout <= #DLY 32'h26486e3e;
				8'h51 : r_dout <= #DLY 32'h8bd78a70;
				8'h52 : r_dout <= #DLY 32'h7477e4c1;
				8'h53 : r_dout <= #DLY 32'hb506e07c;
				8'h54 : r_dout <= #DLY 32'hf32d0a25;
				8'h55 : r_dout <= #DLY 32'h79098b02;
				8'h56 : r_dout <= #DLY 32'he4eabb81;
				8'h57 : r_dout <= #DLY 32'h28123b23;
				8'h58 : r_dout <= #DLY 32'h69dead38;
				8'h59 : r_dout <= #DLY 32'h1574ca16;
				8'h5a : r_dout <= #DLY 32'hdf871b62;
				8'h5b : r_dout <= #DLY 32'h211c40b7;
				8'h5c : r_dout <= #DLY 32'ha51a9ef9;
				8'h5d : r_dout <= #DLY 32'h0014377b;
				8'h5e : r_dout <= #DLY 32'h041e8ac8;
				8'h5f : r_dout <= #DLY 32'h09114003;
				8'h60 : r_dout <= #DLY 32'hbd59e4d2;
				8'h61 : r_dout <= #DLY 32'he3d156d5;
				8'h62 : r_dout <= #DLY 32'h4fe876d5;
				8'h63 : r_dout <= #DLY 32'h2f91a340;
				8'h64 : r_dout <= #DLY 32'h557be8de;
				8'h65 : r_dout <= #DLY 32'h00eae4a7;
				8'h66 : r_dout <= #DLY 32'h0ce5c2ec;
				8'h67 : r_dout <= #DLY 32'h4db4bba6;
				8'h68 : r_dout <= #DLY 32'he756bdff;
				8'h69 : r_dout <= #DLY 32'hdd3369ac;
				8'h6a : r_dout <= #DLY 32'hec17b035;
				8'h6b : r_dout <= #DLY 32'h06572327;
				8'h6c : r_dout <= #DLY 32'h99afc8b0;
				8'h6d : r_dout <= #DLY 32'h56c8c391;
				8'h6e : r_dout <= #DLY 32'h6b65811c;
				8'h6f : r_dout <= #DLY 32'h5e146119;
				8'h70 : r_dout <= #DLY 32'h6e85cb75;
				8'h71 : r_dout <= #DLY 32'hbe07c002;
				8'h72 : r_dout <= #DLY 32'hc2325577;
				8'h73 : r_dout <= #DLY 32'h893ff4ec;
				8'h74 : r_dout <= #DLY 32'h5bbfc92d;
				8'h75 : r_dout <= #DLY 32'hd0ec3b25;
				8'h76 : r_dout <= #DLY 32'hb7801ab7;
				8'h77 : r_dout <= #DLY 32'h8d6d3b24;
				8'h78 : r_dout <= #DLY 32'h20c763ef;
				8'h79 : r_dout <= #DLY 32'hc366a5fc;
				8'h7a : r_dout <= #DLY 32'h9c382880;
				8'h7b : r_dout <= #DLY 32'h0ace3205;
				8'h7c : r_dout <= #DLY 32'haac9548a;
				8'h7d : r_dout <= #DLY 32'heca1d7c7;
				8'h7e : r_dout <= #DLY 32'h041afa32;
				8'h7f : r_dout <= #DLY 32'h1d16625a;
				8'h80 : r_dout <= #DLY 32'h6701902c;
				8'h81 : r_dout <= #DLY 32'h9b757a54;
				8'h82 : r_dout <= #DLY 32'h31d477f7;
				8'h83 : r_dout <= #DLY 32'h9126b031;
				8'h84 : r_dout <= #DLY 32'h36cc6fdb;
				8'h85 : r_dout <= #DLY 32'hc70b8b46;
				8'h86 : r_dout <= #DLY 32'hd9e66a48;
				8'h87 : r_dout <= #DLY 32'h56e55a79;
				8'h88 : r_dout <= #DLY 32'h026a4ceb;
				8'h89 : r_dout <= #DLY 32'h52437eff;
				8'h8a : r_dout <= #DLY 32'h2f8f76b4;
				8'h8b : r_dout <= #DLY 32'h0df980a5;
				8'h8c : r_dout <= #DLY 32'h8674cde3;
				8'h8d : r_dout <= #DLY 32'hedda04eb;
				8'h8e : r_dout <= #DLY 32'h17a9be04;
				8'h8f : r_dout <= #DLY 32'h2c18f4df;
				8'h90 : r_dout <= #DLY 32'hb7747f9d;
				8'h91 : r_dout <= #DLY 32'hab2af7b4;
				8'h92 : r_dout <= #DLY 32'hefc34d20;
				8'h93 : r_dout <= #DLY 32'h2e096b7c;
				8'h94 : r_dout <= #DLY 32'h1741a254;
				8'h95 : r_dout <= #DLY 32'he5b6a035;
				8'h96 : r_dout <= #DLY 32'h213d42f6;
				8'h97 : r_dout <= #DLY 32'h2c1c7c26;
				8'h98 : r_dout <= #DLY 32'h61c2f50f;
				8'h99 : r_dout <= #DLY 32'h6552daf9;
				8'h9a : r_dout <= #DLY 32'hd2c231f8;
				8'h9b : r_dout <= #DLY 32'h25130f69;
				8'h9c : r_dout <= #DLY 32'hd8167fa2;
				8'h9d : r_dout <= #DLY 32'h0418f2c8;
				8'h9e : r_dout <= #DLY 32'h001a96a6;
				8'h9f : r_dout <= #DLY 32'h0d1526ab;
				8'ha0 : r_dout <= #DLY 32'h63315c21;
				8'ha1 : r_dout <= #DLY 32'h5e0a72ec;
				8'ha2 : r_dout <= #DLY 32'h49bafefd;
				8'ha3 : r_dout <= #DLY 32'h187908d9;
				8'ha4 : r_dout <= #DLY 32'h8d0dbd86;
				8'ha5 : r_dout <= #DLY 32'h311170a7;
				8'ha6 : r_dout <= #DLY 32'h3e9b640c;
				8'ha7 : r_dout <= #DLY 32'hcc3e10d7;
				8'ha8 : r_dout <= #DLY 32'hd5cad3b6;
				8'ha9 : r_dout <= #DLY 32'h0caec388;
				8'haa : r_dout <= #DLY 32'hf73001e1;
				8'hab : r_dout <= #DLY 32'h6c728aff;
				8'hac : r_dout <= #DLY 32'h71eae2a1;
				8'had : r_dout <= #DLY 32'h1f9af36e;
				8'hae : r_dout <= #DLY 32'hcfcbd12f;
				8'haf : r_dout <= #DLY 32'hc1de8417;
				8'hb0 : r_dout <= #DLY 32'hac07be6b;
				8'hb1 : r_dout <= #DLY 32'hcb44a1d8;
				8'hb2 : r_dout <= #DLY 32'h8b9b0f56;
				8'hb3 : r_dout <= #DLY 32'h013988c3;
				8'hb4 : r_dout <= #DLY 32'hb1c52fca;
				8'hb5 : r_dout <= #DLY 32'hb4be31cd;
				8'hb6 : r_dout <= #DLY 32'hd8782806;
				8'hb7 : r_dout <= #DLY 32'h12a3a4e2;
				8'hb8 : r_dout <= #DLY 32'h6f7de532;
				8'hb9 : r_dout <= #DLY 32'h58fd7eb6;
				8'hba : r_dout <= #DLY 32'hd01ee900;
				8'hbb : r_dout <= #DLY 32'h24adffc2;
				8'hbc : r_dout <= #DLY 32'hf4990fc5;
				8'hbd : r_dout <= #DLY 32'h9711aac5;
				8'hbe : r_dout <= #DLY 32'h001d7b95;
				8'hbf : r_dout <= #DLY 32'h82e5e7d2;
				8'hc0 : r_dout <= #DLY 32'h109873f6;
				8'hc1 : r_dout <= #DLY 32'h00613096;
				8'hc2 : r_dout <= #DLY 32'hc32d9521;
				8'hc3 : r_dout <= #DLY 32'hada121ff;
				8'hc4 : r_dout <= #DLY 32'h29908415;
				8'hc5 : r_dout <= #DLY 32'h7fbb977f;
				8'hc6 : r_dout <= #DLY 32'haf9eb3db;
				8'hc7 : r_dout <= #DLY 32'h29c9ed2a;
				8'hc8 : r_dout <= #DLY 32'h5ce2a465;
				8'hc9 : r_dout <= #DLY 32'ha730f32c;
				8'hca : r_dout <= #DLY 32'hd0aa3fe8;
				8'hcb : r_dout <= #DLY 32'h8a5cc091;
				8'hcc : r_dout <= #DLY 32'hd49e2ce7;
				8'hcd : r_dout <= #DLY 32'h0ce454a9;
				8'hce : r_dout <= #DLY 32'hd60acd86;
				8'hcf : r_dout <= #DLY 32'h015f1919;
				8'hd0 : r_dout <= #DLY 32'h77079103;
				8'hd1 : r_dout <= #DLY 32'hdea03af6;
				8'hd2 : r_dout <= #DLY 32'h78a8565e;
				8'hd3 : r_dout <= #DLY 32'hdee356df;
				8'hd4 : r_dout <= #DLY 32'h21f05cbe;
				8'hd5 : r_dout <= #DLY 32'h8b75e387;
				8'hd6 : r_dout <= #DLY 32'hb3c50651;
				8'hd7 : r_dout <= #DLY 32'hb8a5c3ef;
				8'hd8 : r_dout <= #DLY 32'hd8eeb6d2;
				8'hd9 : r_dout <= #DLY 32'he523be77;
				8'hda : r_dout <= #DLY 32'hc2154529;
				8'hdb : r_dout <= #DLY 32'h2f69efdf;
				8'hdc : r_dout <= #DLY 32'hafe67afb;
				8'hdd : r_dout <= #DLY 32'hf470c4b2;
				8'hde : r_dout <= #DLY 32'hf3e0eb5b;
				8'hdf : r_dout <= #DLY 32'hd6cc9876;
				8'he0 : r_dout <= #DLY 32'h39e4460c;
				8'he1 : r_dout <= #DLY 32'h1fda8538;
				8'he2 : r_dout <= #DLY 32'h1987832f;
				8'he3 : r_dout <= #DLY 32'hca007367;
				8'he4 : r_dout <= #DLY 32'ha99144f8;
				8'he5 : r_dout <= #DLY 32'h296b299e;
				8'he6 : r_dout <= #DLY 32'h492fc295;
				8'he7 : r_dout <= #DLY 32'h9266beab;
				8'he8 : r_dout <= #DLY 32'hb5676e69;
				8'he9 : r_dout <= #DLY 32'h9bd3ddda;
				8'hea : r_dout <= #DLY 32'hdf7e052f;
				8'heb : r_dout <= #DLY 32'hdb25701c;
				8'hec : r_dout <= #DLY 32'h1b5e51ee;
				8'hed : r_dout <= #DLY 32'hf65324e6;
				8'hee : r_dout <= #DLY 32'h6afce36c;
				8'hef : r_dout <= #DLY 32'h0316cc04;
				8'hf0 : r_dout <= #DLY 32'h8644213e;
				8'hf1 : r_dout <= #DLY 32'hb7dc59d0;
				8'hf2 : r_dout <= #DLY 32'h7965291f;
				8'hf3 : r_dout <= #DLY 32'hccd6fd43;
				8'hf4 : r_dout <= #DLY 32'h41823979;
				8'hf5 : r_dout <= #DLY 32'h932bcdf6;
				8'hf6 : r_dout <= #DLY 32'hb657c34d;
				8'hf7 : r_dout <= #DLY 32'h4edfd282;
				8'hf8 : r_dout <= #DLY 32'h7ae5290c;
				8'hf9 : r_dout <= #DLY 32'h3cb9536b;
				8'hfa : r_dout <= #DLY 32'h851e20fe;
				8'hfb : r_dout <= #DLY 32'h9833557e;
				8'hfc : r_dout <= #DLY 32'h13ecf0b0;
				8'hfd : r_dout <= #DLY 32'hd3ffb372;
				8'hfe : r_dout <= #DLY 32'h3f85c5c1;
				8'hff : r_dout <= #DLY 32'h0aef7ed2;
			endcase
		end else begin
			case(i_addr)  //s-box8
				8'h00 : r_dout <= #DLY 32'he216300d;
				8'h01 : r_dout <= #DLY 32'hbbddfffc;
				8'h02 : r_dout <= #DLY 32'ha7ebdabd;
				8'h03 : r_dout <= #DLY 32'h35648095;
				8'h04 : r_dout <= #DLY 32'h7789f8b7;
				8'h05 : r_dout <= #DLY 32'he6c1121b;
				8'h06 : r_dout <= #DLY 32'h0e241600;
				8'h07 : r_dout <= #DLY 32'h052ce8b5;
				8'h08 : r_dout <= #DLY 32'h11a9cfb0;
				8'h09 : r_dout <= #DLY 32'he5952f11;
				8'h0a : r_dout <= #DLY 32'hece7990a;
				8'h0b : r_dout <= #DLY 32'h9386d174;
				8'h0c : r_dout <= #DLY 32'h2a42931c;
				8'h0d : r_dout <= #DLY 32'h76e38111;
				8'h0e : r_dout <= #DLY 32'hb12def3a;
				8'h0f : r_dout <= #DLY 32'h37ddddfc;
				8'h10 : r_dout <= #DLY 32'hde9adeb1;
				8'h11 : r_dout <= #DLY 32'h0a0cc32c;
				8'h12 : r_dout <= #DLY 32'hbe197029;
				8'h13 : r_dout <= #DLY 32'h84a00940;
				8'h14 : r_dout <= #DLY 32'hbb243a0f;
				8'h15 : r_dout <= #DLY 32'hb4d137cf;
				8'h16 : r_dout <= #DLY 32'hb44e79f0;
				8'h17 : r_dout <= #DLY 32'h049eedfd;
				8'h18 : r_dout <= #DLY 32'h0b15a15d;
				8'h19 : r_dout <= #DLY 32'h480d3168;
				8'h1a : r_dout <= #DLY 32'h8bbbde5a;
				8'h1b : r_dout <= #DLY 32'h669ded42;
				8'h1c : r_dout <= #DLY 32'hc7ece831;
				8'h1d : r_dout <= #DLY 32'h3f8f95e7;
				8'h1e : r_dout <= #DLY 32'h72df191b;
				8'h1f : r_dout <= #DLY 32'h7580330d;
				8'h20 : r_dout <= #DLY 32'h94074251;
				8'h21 : r_dout <= #DLY 32'h5c7dcdfa;
				8'h22 : r_dout <= #DLY 32'habbe6d63;
				8'h23 : r_dout <= #DLY 32'haa402164;
				8'h24 : r_dout <= #DLY 32'hb301d40a;
				8'h25 : r_dout <= #DLY 32'h02e7d1ca;
				8'h26 : r_dout <= #DLY 32'h53571dae;
				8'h27 : r_dout <= #DLY 32'h7a3182a2;
				8'h28 : r_dout <= #DLY 32'h12a8ddec;
				8'h29 : r_dout <= #DLY 32'hfdaa335d;
				8'h2a : r_dout <= #DLY 32'h176f43e8;
				8'h2b : r_dout <= #DLY 32'h71fb46d4;
				8'h2c : r_dout <= #DLY 32'h38129022;
				8'h2d : r_dout <= #DLY 32'hce949ad4;
				8'h2e : r_dout <= #DLY 32'hb84769ad;
				8'h2f : r_dout <= #DLY 32'h965bd862;
				8'h30 : r_dout <= #DLY 32'h82f3d055;
				8'h31 : r_dout <= #DLY 32'h66fb9767;
				8'h32 : r_dout <= #DLY 32'h15b80b4e;
				8'h33 : r_dout <= #DLY 32'h1d5b47a0;
				8'h34 : r_dout <= #DLY 32'h4cfde06f;
				8'h35 : r_dout <= #DLY 32'hc28ec4b8;
				8'h36 : r_dout <= #DLY 32'h57e8726e;
				8'h37 : r_dout <= #DLY 32'h647a78fc;
				8'h38 : r_dout <= #DLY 32'h99865d44;
				8'h39 : r_dout <= #DLY 32'h608bd593;
				8'h3a : r_dout <= #DLY 32'h6c200e03;
				8'h3b : r_dout <= #DLY 32'h39dc5ff6;
				8'h3c : r_dout <= #DLY 32'h5d0b00a3;
				8'h3d : r_dout <= #DLY 32'hae63aff2;
				8'h3e : r_dout <= #DLY 32'h7e8bd632;
				8'h3f : r_dout <= #DLY 32'h70108c0c;
				8'h40 : r_dout <= #DLY 32'hbbd35049;
				8'h41 : r_dout <= #DLY 32'h2998df04;
				8'h42 : r_dout <= #DLY 32'h980cf42a;
				8'h43 : r_dout <= #DLY 32'h9b6df491;
				8'h44 : r_dout <= #DLY 32'h9e7edd53;
				8'h45 : r_dout <= #DLY 32'h06918548;
				8'h46 : r_dout <= #DLY 32'h58cb7e07;
				8'h47 : r_dout <= #DLY 32'h3b74ef2e;
				8'h48 : r_dout <= #DLY 32'h522fffb1;
				8'h49 : r_dout <= #DLY 32'hd24708cc;
				8'h4a : r_dout <= #DLY 32'h1c7e27cd;
				8'h4b : r_dout <= #DLY 32'ha4eb215b;
				8'h4c : r_dout <= #DLY 32'h3cf1d2e2;
				8'h4d : r_dout <= #DLY 32'h19b47a38;
				8'h4e : r_dout <= #DLY 32'h424f7618;
				8'h4f : r_dout <= #DLY 32'h35856039;
				8'h50 : r_dout <= #DLY 32'h9d17dee7;
				8'h51 : r_dout <= #DLY 32'h27eb35e6;
				8'h52 : r_dout <= #DLY 32'hc9aff67b;
				8'h53 : r_dout <= #DLY 32'h36baf5b8;
				8'h54 : r_dout <= #DLY 32'h09c467cd;
				8'h55 : r_dout <= #DLY 32'hc18910b1;
				8'h56 : r_dout <= #DLY 32'he11dbf7b;
				8'h57 : r_dout <= #DLY 32'h06cd1af8;
				8'h58 : r_dout <= #DLY 32'h7170c608;
				8'h59 : r_dout <= #DLY 32'h2d5e3354;
				8'h5a : r_dout <= #DLY 32'hd4de495a;
				8'h5b : r_dout <= #DLY 32'h64c6d006;
				8'h5c : r_dout <= #DLY 32'hbcc0c62c;
				8'h5d : r_dout <= #DLY 32'h3dd00db3;
				8'h5e : r_dout <= #DLY 32'h708f8f34;
				8'h5f : r_dout <= #DLY 32'h77d51b42;
				8'h60 : r_dout <= #DLY 32'h264f620f;
				8'h61 : r_dout <= #DLY 32'h24b8d2bf;
				8'h62 : r_dout <= #DLY 32'h15c1b79e;
				8'h63 : r_dout <= #DLY 32'h46a52564;
				8'h64 : r_dout <= #DLY 32'hf8d7e54e;
				8'h65 : r_dout <= #DLY 32'h3e378160;
				8'h66 : r_dout <= #DLY 32'h7895cda5;
				8'h67 : r_dout <= #DLY 32'h859c15a5;
				8'h68 : r_dout <= #DLY 32'he6459788;
				8'h69 : r_dout <= #DLY 32'hc37bc75f;
				8'h6a : r_dout <= #DLY 32'hdb07ba0c;
				8'h6b : r_dout <= #DLY 32'h0676a3ab;
				8'h6c : r_dout <= #DLY 32'h7f229b1e;
				8'h6d : r_dout <= #DLY 32'h31842e7b;
				8'h6e : r_dout <= #DLY 32'h24259fd7;
				8'h6f : r_dout <= #DLY 32'hf8bef472;
				8'h70 : r_dout <= #DLY 32'h835ffcb8;
				8'h71 : r_dout <= #DLY 32'h6df4c1f2;
				8'h72 : r_dout <= #DLY 32'h96f5b195;
				8'h73 : r_dout <= #DLY 32'hfd0af0fc;
				8'h74 : r_dout <= #DLY 32'hb0fe134c;
				8'h75 : r_dout <= #DLY 32'he2506d3d;
				8'h76 : r_dout <= #DLY 32'h4f9b12ea;
				8'h77 : r_dout <= #DLY 32'hf215f225;
				8'h78 : r_dout <= #DLY 32'ha223736f;
				8'h79 : r_dout <= #DLY 32'h9fb4c428;
				8'h7a : r_dout <= #DLY 32'h25d04979;
				8'h7b : r_dout <= #DLY 32'h34c713f8;
				8'h7c : r_dout <= #DLY 32'hc4618187;
				8'h7d : r_dout <= #DLY 32'hea7a6e98;
				8'h7e : r_dout <= #DLY 32'h7cd16efc;
				8'h7f : r_dout <= #DLY 32'h1436876c;
				8'h80 : r_dout <= #DLY 32'hf1544107;
				8'h81 : r_dout <= #DLY 32'hbedeee14;
				8'h82 : r_dout <= #DLY 32'h56e9af27;
				8'h83 : r_dout <= #DLY 32'ha04aa441;
				8'h84 : r_dout <= #DLY 32'h3cf7c899;
				8'h85 : r_dout <= #DLY 32'h92ecbae6;
				8'h86 : r_dout <= #DLY 32'hdd67016d;
				8'h87 : r_dout <= #DLY 32'h151682eb;
				8'h88 : r_dout <= #DLY 32'ha842eedf;
				8'h89 : r_dout <= #DLY 32'hfdba60b4;
				8'h8a : r_dout <= #DLY 32'hf1907b75;
				8'h8b : r_dout <= #DLY 32'h20e3030f;
				8'h8c : r_dout <= #DLY 32'h24d8c29e;
				8'h8d : r_dout <= #DLY 32'he139673b;
				8'h8e : r_dout <= #DLY 32'hefa63fb8;
				8'h8f : r_dout <= #DLY 32'h71873054;
				8'h90 : r_dout <= #DLY 32'hb6f2cf3b;
				8'h91 : r_dout <= #DLY 32'h9f326442;
				8'h92 : r_dout <= #DLY 32'hcb15a4cc;
				8'h93 : r_dout <= #DLY 32'hb01a4504;
				8'h94 : r_dout <= #DLY 32'hf1e47d8d;
				8'h95 : r_dout <= #DLY 32'h844a1be5;
				8'h96 : r_dout <= #DLY 32'hbae7dfdc;
				8'h97 : r_dout <= #DLY 32'h42cbda70;
				8'h98 : r_dout <= #DLY 32'hcd7dae0a;
				8'h99 : r_dout <= #DLY 32'h57e85b7a;
				8'h9a : r_dout <= #DLY 32'hd53f5af6;
				8'h9b : r_dout <= #DLY 32'h20cf4d8c;
				8'h9c : r_dout <= #DLY 32'hcea4d428;
				8'h9d : r_dout <= #DLY 32'h79d130a4;
				8'h9e : r_dout <= #DLY 32'h3486ebfb;
				8'h9f : r_dout <= #DLY 32'h33d3cddc;
				8'ha0 : r_dout <= #DLY 32'h77853b53;
				8'ha1 : r_dout <= #DLY 32'h37effcb5;
				8'ha2 : r_dout <= #DLY 32'hc5068778;
				8'ha3 : r_dout <= #DLY 32'he580b3e6;
				8'ha4 : r_dout <= #DLY 32'h4e68b8f4;
				8'ha5 : r_dout <= #DLY 32'hc5c8b37e;
				8'ha6 : r_dout <= #DLY 32'h0d809ea2;
				8'ha7 : r_dout <= #DLY 32'h398feb7c;
				8'ha8 : r_dout <= #DLY 32'h132a4f94;
				8'ha9 : r_dout <= #DLY 32'h43b7950e;
				8'haa : r_dout <= #DLY 32'h2fee7d1c;
				8'hab : r_dout <= #DLY 32'h223613bd;
				8'hac : r_dout <= #DLY 32'hdd06caa2;
				8'had : r_dout <= #DLY 32'h37df932b;
				8'hae : r_dout <= #DLY 32'hc4248289;
				8'haf : r_dout <= #DLY 32'hacf3ebc3;
				8'hb0 : r_dout <= #DLY 32'h5715f6b7;
				8'hb1 : r_dout <= #DLY 32'hef3478dd;
				8'hb2 : r_dout <= #DLY 32'hf267616f;
				8'hb3 : r_dout <= #DLY 32'hc148cbe4;
				8'hb4 : r_dout <= #DLY 32'h9052815e;
				8'hb5 : r_dout <= #DLY 32'h5e410fab;
				8'hb6 : r_dout <= #DLY 32'hb48a2465;
				8'hb7 : r_dout <= #DLY 32'h2eda7fa4;
				8'hb8 : r_dout <= #DLY 32'he87b40e4;
				8'hb9 : r_dout <= #DLY 32'he98ea084;
				8'hba : r_dout <= #DLY 32'h5889e9e1;
				8'hbb : r_dout <= #DLY 32'hefd390fc;
				8'hbc : r_dout <= #DLY 32'hdd07d35b;
				8'hbd : r_dout <= #DLY 32'hdb485694;
				8'hbe : r_dout <= #DLY 32'h38d7e5b2;
				8'hbf : r_dout <= #DLY 32'h57720101;
				8'hc0 : r_dout <= #DLY 32'h730edebc;
				8'hc1 : r_dout <= #DLY 32'h5b643113;
				8'hc2 : r_dout <= #DLY 32'h94917e4f;
				8'hc3 : r_dout <= #DLY 32'h503c2fba;
				8'hc4 : r_dout <= #DLY 32'h646f1282;
				8'hc5 : r_dout <= #DLY 32'h7523d24a;
				8'hc6 : r_dout <= #DLY 32'he0779695;
				8'hc7 : r_dout <= #DLY 32'hf9c17a8f;
				8'hc8 : r_dout <= #DLY 32'h7a5b2121;
				8'hc9 : r_dout <= #DLY 32'hd187b896;
				8'hca : r_dout <= #DLY 32'h29263a4d;
				8'hcb : r_dout <= #DLY 32'hba510cdf;
				8'hcc : r_dout <= #DLY 32'h81f47c9f;
				8'hcd : r_dout <= #DLY 32'had1163ed;
				8'hce : r_dout <= #DLY 32'hea7b5965;
				8'hcf : r_dout <= #DLY 32'h1a00726e;
				8'hd0 : r_dout <= #DLY 32'h11403092;
				8'hd1 : r_dout <= #DLY 32'h00da6d77;
				8'hd2 : r_dout <= #DLY 32'h4a0cdd61;
				8'hd3 : r_dout <= #DLY 32'had1f4603;
				8'hd4 : r_dout <= #DLY 32'h605bdfb0;
				8'hd5 : r_dout <= #DLY 32'h9eedc364;
				8'hd6 : r_dout <= #DLY 32'h22ebe6a8;
				8'hd7 : r_dout <= #DLY 32'hcee7d28a;
				8'hd8 : r_dout <= #DLY 32'ha0e736a0;
				8'hd9 : r_dout <= #DLY 32'h5564a6b9;
				8'hda : r_dout <= #DLY 32'h10853209;
				8'hdb : r_dout <= #DLY 32'hc7eb8f37;
				8'hdc : r_dout <= #DLY 32'h2de705ca;
				8'hdd : r_dout <= #DLY 32'h8951570f;
				8'hde : r_dout <= #DLY 32'hdf09822b;
				8'hdf : r_dout <= #DLY 32'hbd691a6c;
				8'he0 : r_dout <= #DLY 32'haa12e4f2;
				8'he1 : r_dout <= #DLY 32'h87451c0f;
				8'he2 : r_dout <= #DLY 32'he0f6a27a;
				8'he3 : r_dout <= #DLY 32'h3ada4819;
				8'he4 : r_dout <= #DLY 32'h4cf1764f;
				8'he5 : r_dout <= #DLY 32'h0d771c2b;
				8'he6 : r_dout <= #DLY 32'h67cdb156;
				8'he7 : r_dout <= #DLY 32'h350d8384;
				8'he8 : r_dout <= #DLY 32'h5938fa0f;
				8'he9 : r_dout <= #DLY 32'h42399ef3;
				8'hea : r_dout <= #DLY 32'h36997b07;
				8'heb : r_dout <= #DLY 32'h0e84093d;
				8'hec : r_dout <= #DLY 32'h4aa93e61;
				8'hed : r_dout <= #DLY 32'h8360d87b;
				8'hee : r_dout <= #DLY 32'h1fa98b0c;
				8'hef : r_dout <= #DLY 32'h1149382c;
				8'hf0 : r_dout <= #DLY 32'he97625a5;
				8'hf1 : r_dout <= #DLY 32'h0614d1b7;
				8'hf2 : r_dout <= #DLY 32'h0e25244b;
				8'hf3 : r_dout <= #DLY 32'h0c768347;
				8'hf4 : r_dout <= #DLY 32'h589e8d82;
				8'hf5 : r_dout <= #DLY 32'h0d2059d1;
				8'hf6 : r_dout <= #DLY 32'ha466bb1e;
				8'hf7 : r_dout <= #DLY 32'hf8da0a82;
				8'hf8 : r_dout <= #DLY 32'h04f19130;
				8'hf9 : r_dout <= #DLY 32'hba6e4ec0;
				8'hfa : r_dout <= #DLY 32'h99265164;
				8'hfb : r_dout <= #DLY 32'h1ee7230d;
				8'hfc : r_dout <= #DLY 32'h50b2ad80;
				8'hfd : r_dout <= #DLY 32'heaee6801;
				8'hfe : r_dout <= #DLY 32'h8db2a283;
				8'hff : r_dout <= #DLY 32'hea8bf59e;
			endcase
		end		
    end

endmodule
